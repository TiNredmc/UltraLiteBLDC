-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 20 2022 14:33:48

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    LED_G : out std_logic;
    io_i2c_sda : inout std_logic;
    io_i2c_scl : in std_logic;
    LED_R : out std_logic;
    LED_B : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2565\ : std_logic;
signal \N__2562\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2532\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2487\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2388\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2337\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2307\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2247\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2211\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2180\ : std_logic;
signal \N__2177\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2162\ : std_logic;
signal \N__2159\ : std_logic;
signal \N__2154\ : std_logic;
signal \N__2151\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2145\ : std_logic;
signal \N__2142\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2136\ : std_logic;
signal \N__2133\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2127\ : std_logic;
signal \N__2124\ : std_logic;
signal \N__2121\ : std_logic;
signal \N__2118\ : std_logic;
signal \N__2115\ : std_logic;
signal \N__2112\ : std_logic;
signal \N__2109\ : std_logic;
signal \N__2106\ : std_logic;
signal \N__2103\ : std_logic;
signal \N__2100\ : std_logic;
signal \N__2097\ : std_logic;
signal \N__2094\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2088\ : std_logic;
signal \N__2085\ : std_logic;
signal \N__2082\ : std_logic;
signal \N__2079\ : std_logic;
signal \N__2076\ : std_logic;
signal \N__2073\ : std_logic;
signal \N__2070\ : std_logic;
signal \N__2067\ : std_logic;
signal \N__2064\ : std_logic;
signal \N__2061\ : std_logic;
signal \N__2058\ : std_logic;
signal \N__2055\ : std_logic;
signal \N__2052\ : std_logic;
signal \N__2049\ : std_logic;
signal \N__2046\ : std_logic;
signal \N__2043\ : std_logic;
signal \N__2040\ : std_logic;
signal \N__2037\ : std_logic;
signal \N__2034\ : std_logic;
signal \N__2031\ : std_logic;
signal \N__2028\ : std_logic;
signal \N__2025\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal sdaoe_i : std_logic;
signal sdaout_i : std_logic;
signal sdain_i : std_logic;
signal sclin_i : std_logic;
signal \n2965_cascade_\ : std_logic;
signal \n2870_cascade_\ : std_logic;
signal \n6_adj_16_cascade_\ : std_logic;
signal n2967 : std_logic;
signal n2966 : std_logic;
signal \n2811_cascade_\ : std_logic;
signal \n2821_cascade_\ : std_logic;
signal \n1_adj_12_cascade_\ : std_logic;
signal \PWM_B\ : std_logic;
signal \PWM_G\ : std_logic;
signal \PWM_R\ : std_logic;
signal n1815 : std_logic;
signal n1_adj_12 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \hard0_SBDATo_0\ : std_logic;
signal \hard0_SBDATo_1\ : std_logic;
signal \hard0_SBDATo_3\ : std_logic;
signal \hard0_SBDATo_4\ : std_logic;
signal \hard0_SBDATo_5\ : std_logic;
signal \hard0_SBDATo_7\ : std_logic;
signal i2c_cmd_1_0 : std_logic;
signal i2c_cmd_1_1 : std_logic;
signal i2c_cmd_1_2 : std_logic;
signal \PWM_duty_2\ : std_logic;
signal i2c_cmd_1_5 : std_logic;
signal i2c_cmd_1_6 : std_logic;
signal i2c_cmd_1_7 : std_logic;
signal i2c_cmd_1_4 : std_logic;
signal i2c_cmd_1_3 : std_logic;
signal \bfn_1_4_0_\ : std_logic;
signal n2514 : std_logic;
signal n2515 : std_logic;
signal n2516 : std_logic;
signal n2517 : std_logic;
signal n2518 : std_logic;
signal n2519 : std_logic;
signal n2520 : std_logic;
signal n1831 : std_logic;
signal \n12_adj_11_cascade_\ : std_logic;
signal n4_adj_15 : std_logic;
signal n8 : std_logic;
signal \n14_cascade_\ : std_logic;
signal n2012 : std_logic;
signal n2955 : std_logic;
signal drv_cnt_1 : std_logic;
signal drv_cnt_0 : std_logic;
signal \n2955_cascade_\ : std_logic;
signal drv_cnt_2 : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal n2521 : std_logic;
signal n2522 : std_logic;
signal n2523 : std_logic;
signal n2524 : std_logic;
signal n2525 : std_logic;
signal drv_clk_counter_6 : std_logic;
signal n2526 : std_logic;
signal drv_clk_counter_7 : std_logic;
signal n2527 : std_logic;
signal n2528 : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal n2529 : std_logic;
signal n2530 : std_logic;
signal \n2838_cascade_\ : std_logic;
signal i2c_cmd_0_5 : std_logic;
signal i2c_cmd_0_6 : std_logic;
signal i2c_cmd_0_3 : std_logic;
signal \n6_adj_8_cascade_\ : std_logic;
signal i2c_cmd_0_7 : std_logic;
signal i2c_cmd_0_2 : std_logic;
signal n10_adj_2 : std_logic;
signal \n17_adj_18_cascade_\ : std_logic;
signal \PWM_cnt_2\ : std_logic;
signal \PWM_cnt_3\ : std_logic;
signal \PWM_duty_3\ : std_logic;
signal \PWM_duty_4\ : std_logic;
signal \n6_adj_5_cascade_\ : std_logic;
signal \PWM_cnt_4\ : std_logic;
signal n2247 : std_logic;
signal \n2250_cascade_\ : std_logic;
signal i2c_cmd_0_1 : std_logic;
signal i2c_cmd_0_4 : std_logic;
signal i2c_cmd_0_0 : std_logic;
signal n2858 : std_logic;
signal n1778 : std_logic;
signal \PWM_duty_5\ : std_logic;
signal n2968 : std_logic;
signal n2883 : std_logic;
signal \n2883_cascade_\ : std_logic;
signal \PWM_duty_0\ : std_logic;
signal \PWM_cnt_1\ : std_logic;
signal \PWM_cnt_0\ : std_logic;
signal \PWM_duty_1\ : std_logic;
signal n4_adj_17 : std_logic;
signal \PWM_duty_6\ : std_logic;
signal \PWM_cnt_6\ : std_logic;
signal \PWM_cnt_5\ : std_logic;
signal \n10_cascade_\ : std_logic;
signal n12_adj_13 : std_logic;
signal n8_adj_10 : std_logic;
signal n2881 : std_logic;
signal n14_adj_14 : std_logic;
signal \n104_cascade_\ : std_logic;
signal n105 : std_logic;
signal n1921 : std_logic;
signal \PWM_duty_7\ : std_logic;
signal \PWM_cnt_7\ : std_logic;
signal n2969 : std_logic;
signal drv_clk_counter_4 : std_logic;
signal drv_clk_counter_1 : std_logic;
signal drv_clk_counter_0 : std_logic;
signal drv_clk_counter_8 : std_logic;
signal drv_clk_counter_5 : std_logic;
signal \n2810_cascade_\ : std_logic;
signal n2819 : std_logic;
signal motor_on : std_logic;
signal drv_clk_counter_10 : std_logic;
signal \n2820_cascade_\ : std_logic;
signal drv_clk_counter_9 : std_logic;
signal n953 : std_logic;
signal drv_clk_counter_2 : std_logic;
signal drv_clk_counter_3 : std_logic;
signal n2963 : std_logic;
signal \n2824_cascade_\ : std_logic;
signal \hard_SBADRi_3\ : std_logic;
signal n2981 : std_logic;
signal \GB_BUFFER_n2981_THRU_CO\ : std_logic;
signal \n2960_cascade_\ : std_logic;
signal \hard_SBWRi\ : std_logic;
signal \hard_SBADRi_0\ : std_logic;
signal \n12_adj_7_cascade_\ : std_logic;
signal \hard_SBADRi_2\ : std_logic;
signal n2971 : std_logic;
signal \n13_adj_6_cascade_\ : std_logic;
signal \hard_SBDATi_4\ : std_logic;
signal \n12_cascade_\ : std_logic;
signal \hard_SBDATi_2\ : std_logic;
signal n15 : std_logic;
signal \n2974_cascade_\ : std_logic;
signal \n2970_cascade_\ : std_logic;
signal \hard_SBSTBi\ : std_logic;
signal n31 : std_logic;
signal n2970 : std_logic;
signal n2243 : std_logic;
signal \n17_cascade_\ : std_logic;
signal \n1887_cascade_\ : std_logic;
signal n1852 : std_logic;
signal n22_adj_9 : std_logic;
signal n2959 : std_logic;
signal n1887 : std_logic;
signal n4 : std_logic;
signal n1779 : std_logic;
signal n2972 : std_logic;
signal \n13_cascade_\ : std_logic;
signal \n4_adj_19_cascade_\ : std_logic;
signal \hard_SBADRi_1\ : std_logic;
signal \n13_adj_4_cascade_\ : std_logic;
signal \hard_SBDATi_7\ : std_logic;
signal cmd_decoded : std_logic;
signal \n2961_cascade_\ : std_logic;
signal n2961 : std_logic;
signal n2973 : std_logic;
signal n2962 : std_logic;
signal \hard0_SBDATo_6\ : std_logic;
signal \i2c_stat_7_N_205_6_cascade_\ : std_logic;
signal i2c_stat_6 : std_logic;
signal i2c_cnt_1 : std_logic;
signal i2c_cnt_0 : std_logic;
signal \n2534_cascade_\ : std_logic;
signal \n25_cascade_\ : std_logic;
signal \hard0_SBDATo_2\ : std_logic;
signal n2534 : std_logic;
signal n4_adj_1 : std_logic;
signal \n2840_cascade_\ : std_logic;
signal n2850 : std_logic;
signal \n29_cascade_\ : std_logic;
signal n26 : std_logic;
signal n2958 : std_logic;
signal \i2c_stat_7_N_205_2\ : std_logic;
signal \n2958_cascade_\ : std_logic;
signal n20 : std_logic;
signal i2c_stat_2 : std_logic;
signal n2964 : std_logic;
signal \hard0_SBACKo\ : std_logic;
signal i2c_steps_1 : std_logic;
signal i2c_steps_2 : std_logic;
signal i2c_steps_0 : std_logic;
signal \n2957_cascade_\ : std_logic;
signal i2c_steps_3 : std_logic;
signal n1780 : std_logic;
signal n1730 : std_logic;
signal i2c_cmd_cnt_1 : std_logic;
signal i2c_cmd_cnt_0 : std_logic;
signal i2c_cmd_cnt_2 : std_logic;
signal \_gnd_net_\ : std_logic;
signal sysclk : std_logic;
signal n2956 : std_logic;
signal n2016 : std_logic;

signal io_i2c_scl_wire : std_logic;
signal \LED_B_wire\ : std_logic;
signal \LED_G_wire\ : std_logic;
signal \LED_R_wire\ : std_logic;

begin
    io_i2c_scl_wire <= io_i2c_scl;
    LED_B <= \LED_B_wire\;
    LED_G <= \LED_G_wire\;
    LED_R <= \LED_R_wire\;

    \sbio_sda_iopad_od\ : IO_PAD_OD
    port map (
            OE => \N__4990\,
            DIN => \N__4989\,
            DOUT => \N__4988\,
            PACKAGEPIN => io_i2c_sda
        );

    \sbio_sda_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4990\,
            PADOUT => \N__4989\,
            PADIN => \N__4988\,
            CLOCKENABLE => 'H',
            DIN0 => sdain_i,
            DOUT0 => \N__2046\,
            OUTPUTCLK => '0',
            DIN1 => OPEN,
            DOUT1 => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTENABLE => \N__2070\,
            INPUTCLK => '0'
        );

    \sbio_scl_iopad_od\ : IO_PAD_OD
    port map (
            OE => \N__4981\,
            DIN => \N__4980\,
            DOUT => \N__4979\,
            PACKAGEPIN => io_i2c_scl_wire
        );

    \sbio_scl_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4981\,
            PADOUT => \N__4980\,
            PADIN => \N__4979\,
            CLOCKENABLE => 'H',
            DIN0 => sclin_i,
            DOUT0 => \GNDG0\,
            OUTPUTCLK => '0',
            DIN1 => OPEN,
            DOUT1 => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTENABLE => '0',
            INPUTCLK => '0'
        );

    \I__1148\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4954\
        );

    \I__1147\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4954\
        );

    \I__1146\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4951\
        );

    \I__1145\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4948\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__4954\,
            I => i2c_stat_2
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__4951\,
            I => i2c_stat_2
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__4948\,
            I => i2c_stat_2
        );

    \I__1141\ : InMux
    port map (
            O => \N__4941\,
            I => \N__4938\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__4938\,
            I => n2964
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__4935\,
            I => \N__4923\
        );

    \I__1138\ : InMux
    port map (
            O => \N__4934\,
            I => \N__4919\
        );

    \I__1137\ : InMux
    port map (
            O => \N__4933\,
            I => \N__4914\
        );

    \I__1136\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4914\
        );

    \I__1135\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4911\
        );

    \I__1134\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4908\
        );

    \I__1133\ : InMux
    port map (
            O => \N__4929\,
            I => \N__4903\
        );

    \I__1132\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4903\
        );

    \I__1131\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4900\
        );

    \I__1130\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4893\
        );

    \I__1129\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4893\
        );

    \I__1128\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4893\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__4919\,
            I => \N__4884\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__4914\,
            I => \N__4884\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__4911\,
            I => \N__4884\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__4908\,
            I => \N__4884\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__4903\,
            I => \N__4872\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__4900\,
            I => \N__4872\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__4893\,
            I => \N__4872\
        );

    \I__1120\ : Span4Mux_s2_v
    port map (
            O => \N__4884\,
            I => \N__4869\
        );

    \I__1119\ : InMux
    port map (
            O => \N__4883\,
            I => \N__4860\
        );

    \I__1118\ : InMux
    port map (
            O => \N__4882\,
            I => \N__4860\
        );

    \I__1117\ : InMux
    port map (
            O => \N__4881\,
            I => \N__4860\
        );

    \I__1116\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4860\
        );

    \I__1115\ : InMux
    port map (
            O => \N__4879\,
            I => \N__4857\
        );

    \I__1114\ : Span12Mux_s2_v
    port map (
            O => \N__4872\,
            I => \N__4848\
        );

    \I__1113\ : Sp12to4
    port map (
            O => \N__4869\,
            I => \N__4848\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__4860\,
            I => \N__4848\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__4857\,
            I => \N__4848\
        );

    \I__1110\ : Odrv12
    port map (
            O => \N__4848\,
            I => \N__4845\
        );

    \I__1109\ : DummyBuf
    port map (
            O => \N__4845\,
            I => \hard0_SBACKo\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__4842\,
            I => \N__4836\
        );

    \I__1107\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4822\
        );

    \I__1106\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4817\
        );

    \I__1105\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4817\
        );

    \I__1104\ : InMux
    port map (
            O => \N__4836\,
            I => \N__4812\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__4835\,
            I => \N__4805\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__4834\,
            I => \N__4802\
        );

    \I__1101\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4792\
        );

    \I__1100\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4792\
        );

    \I__1099\ : InMux
    port map (
            O => \N__4831\,
            I => \N__4792\
        );

    \I__1098\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4789\
        );

    \I__1097\ : InMux
    port map (
            O => \N__4829\,
            I => \N__4784\
        );

    \I__1096\ : InMux
    port map (
            O => \N__4828\,
            I => \N__4784\
        );

    \I__1095\ : InMux
    port map (
            O => \N__4827\,
            I => \N__4779\
        );

    \I__1094\ : InMux
    port map (
            O => \N__4826\,
            I => \N__4779\
        );

    \I__1093\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4776\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__4822\,
            I => \N__4771\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__4817\,
            I => \N__4771\
        );

    \I__1090\ : InMux
    port map (
            O => \N__4816\,
            I => \N__4766\
        );

    \I__1089\ : InMux
    port map (
            O => \N__4815\,
            I => \N__4766\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__4812\,
            I => \N__4763\
        );

    \I__1087\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4760\
        );

    \I__1086\ : InMux
    port map (
            O => \N__4810\,
            I => \N__4753\
        );

    \I__1085\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4753\
        );

    \I__1084\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4753\
        );

    \I__1083\ : InMux
    port map (
            O => \N__4805\,
            I => \N__4742\
        );

    \I__1082\ : InMux
    port map (
            O => \N__4802\,
            I => \N__4742\
        );

    \I__1081\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4742\
        );

    \I__1080\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4742\
        );

    \I__1079\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4742\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__4792\,
            I => i2c_steps_1
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__4789\,
            I => i2c_steps_1
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__4784\,
            I => i2c_steps_1
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__4779\,
            I => i2c_steps_1
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__4776\,
            I => i2c_steps_1
        );

    \I__1073\ : Odrv4
    port map (
            O => \N__4771\,
            I => i2c_steps_1
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__4766\,
            I => i2c_steps_1
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__4763\,
            I => i2c_steps_1
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__4760\,
            I => i2c_steps_1
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__4753\,
            I => i2c_steps_1
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__4742\,
            I => i2c_steps_1
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__4719\,
            I => \N__4704\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__4718\,
            I => \N__4697\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__4717\,
            I => \N__4693\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__4716\,
            I => \N__4690\
        );

    \I__1063\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4685\
        );

    \I__1062\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4685\
        );

    \I__1061\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4676\
        );

    \I__1060\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4676\
        );

    \I__1059\ : InMux
    port map (
            O => \N__4711\,
            I => \N__4676\
        );

    \I__1058\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4676\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__4709\,
            I => \N__4673\
        );

    \I__1056\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4665\
        );

    \I__1055\ : InMux
    port map (
            O => \N__4707\,
            I => \N__4658\
        );

    \I__1054\ : InMux
    port map (
            O => \N__4704\,
            I => \N__4658\
        );

    \I__1053\ : InMux
    port map (
            O => \N__4703\,
            I => \N__4658\
        );

    \I__1052\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4651\
        );

    \I__1051\ : InMux
    port map (
            O => \N__4701\,
            I => \N__4651\
        );

    \I__1050\ : InMux
    port map (
            O => \N__4700\,
            I => \N__4651\
        );

    \I__1049\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4648\
        );

    \I__1048\ : InMux
    port map (
            O => \N__4696\,
            I => \N__4645\
        );

    \I__1047\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4640\
        );

    \I__1046\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4640\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__4685\,
            I => \N__4637\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__4676\,
            I => \N__4634\
        );

    \I__1043\ : InMux
    port map (
            O => \N__4673\,
            I => \N__4631\
        );

    \I__1042\ : InMux
    port map (
            O => \N__4672\,
            I => \N__4626\
        );

    \I__1041\ : InMux
    port map (
            O => \N__4671\,
            I => \N__4626\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4619\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4669\,
            I => \N__4619\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4668\,
            I => \N__4619\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__4665\,
            I => i2c_steps_2
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4658\,
            I => i2c_steps_2
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__4651\,
            I => i2c_steps_2
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__4648\,
            I => i2c_steps_2
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__4645\,
            I => i2c_steps_2
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__4640\,
            I => i2c_steps_2
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__4637\,
            I => i2c_steps_2
        );

    \I__1030\ : Odrv4
    port map (
            O => \N__4634\,
            I => i2c_steps_2
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__4631\,
            I => i2c_steps_2
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4626\,
            I => i2c_steps_2
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__4619\,
            I => i2c_steps_2
        );

    \I__1026\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4591\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4586\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4594\,
            I => \N__4586\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__4591\,
            I => \N__4575\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__4586\,
            I => \N__4572\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4585\,
            I => \N__4565\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4565\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4565\
        );

    \I__1018\ : CascadeMux
    port map (
            O => \N__4582\,
            I => \N__4556\
        );

    \I__1017\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4541\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4580\,
            I => \N__4541\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4541\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4541\
        );

    \I__1013\ : Span4Mux_s1_v
    port map (
            O => \N__4575\,
            I => \N__4534\
        );

    \I__1012\ : Span4Mux_v
    port map (
            O => \N__4572\,
            I => \N__4534\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4565\,
            I => \N__4534\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4564\,
            I => \N__4531\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4563\,
            I => \N__4522\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4562\,
            I => \N__4522\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4561\,
            I => \N__4522\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4522\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4517\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4517\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4510\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4510\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4510\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4503\
        );

    \I__999\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4503\
        );

    \I__998\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4503\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__4541\,
            I => i2c_steps_0
        );

    \I__996\ : Odrv4
    port map (
            O => \N__4534\,
            I => i2c_steps_0
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4531\,
            I => i2c_steps_0
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4522\,
            I => i2c_steps_0
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4517\,
            I => i2c_steps_0
        );

    \I__992\ : LocalMux
    port map (
            O => \N__4510\,
            I => i2c_steps_0
        );

    \I__991\ : LocalMux
    port map (
            O => \N__4503\,
            I => i2c_steps_0
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__4488\,
            I => \n2957_cascade_\
        );

    \I__989\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4467\
        );

    \I__988\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4462\
        );

    \I__987\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4462\
        );

    \I__986\ : InMux
    port map (
            O => \N__4482\,
            I => \N__4459\
        );

    \I__985\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4450\
        );

    \I__984\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4450\
        );

    \I__983\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4450\
        );

    \I__982\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4450\
        );

    \I__981\ : InMux
    port map (
            O => \N__4477\,
            I => \N__4443\
        );

    \I__980\ : InMux
    port map (
            O => \N__4476\,
            I => \N__4443\
        );

    \I__979\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4443\
        );

    \I__978\ : InMux
    port map (
            O => \N__4474\,
            I => \N__4436\
        );

    \I__977\ : InMux
    port map (
            O => \N__4473\,
            I => \N__4436\
        );

    \I__976\ : InMux
    port map (
            O => \N__4472\,
            I => \N__4436\
        );

    \I__975\ : InMux
    port map (
            O => \N__4471\,
            I => \N__4433\
        );

    \I__974\ : InMux
    port map (
            O => \N__4470\,
            I => \N__4430\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4467\,
            I => \N__4427\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4462\,
            I => \N__4418\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4459\,
            I => \N__4418\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4450\,
            I => \N__4411\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4443\,
            I => \N__4411\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__4436\,
            I => \N__4411\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4433\,
            I => \N__4402\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4430\,
            I => \N__4397\
        );

    \I__965\ : Span4Mux_s3_v
    port map (
            O => \N__4427\,
            I => \N__4397\
        );

    \I__964\ : InMux
    port map (
            O => \N__4426\,
            I => \N__4392\
        );

    \I__963\ : InMux
    port map (
            O => \N__4425\,
            I => \N__4392\
        );

    \I__962\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4387\
        );

    \I__961\ : InMux
    port map (
            O => \N__4423\,
            I => \N__4387\
        );

    \I__960\ : Span4Mux_s1_v
    port map (
            O => \N__4418\,
            I => \N__4382\
        );

    \I__959\ : Span4Mux_h
    port map (
            O => \N__4411\,
            I => \N__4382\
        );

    \I__958\ : InMux
    port map (
            O => \N__4410\,
            I => \N__4371\
        );

    \I__957\ : InMux
    port map (
            O => \N__4409\,
            I => \N__4371\
        );

    \I__956\ : InMux
    port map (
            O => \N__4408\,
            I => \N__4371\
        );

    \I__955\ : InMux
    port map (
            O => \N__4407\,
            I => \N__4371\
        );

    \I__954\ : InMux
    port map (
            O => \N__4406\,
            I => \N__4371\
        );

    \I__953\ : InMux
    port map (
            O => \N__4405\,
            I => \N__4368\
        );

    \I__952\ : Odrv4
    port map (
            O => \N__4402\,
            I => i2c_steps_3
        );

    \I__951\ : Odrv4
    port map (
            O => \N__4397\,
            I => i2c_steps_3
        );

    \I__950\ : LocalMux
    port map (
            O => \N__4392\,
            I => i2c_steps_3
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4387\,
            I => i2c_steps_3
        );

    \I__948\ : Odrv4
    port map (
            O => \N__4382\,
            I => i2c_steps_3
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4371\,
            I => i2c_steps_3
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4368\,
            I => i2c_steps_3
        );

    \I__945\ : CEMux
    port map (
            O => \N__4353\,
            I => \N__4350\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4350\,
            I => \N__4347\
        );

    \I__943\ : Span4Mux_s1_v
    port map (
            O => \N__4347\,
            I => \N__4344\
        );

    \I__942\ : Span4Mux_h
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__941\ : Odrv4
    port map (
            O => \N__4341\,
            I => n1780
        );

    \I__940\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__938\ : Span4Mux_s3_h
    port map (
            O => \N__4332\,
            I => \N__4329\
        );

    \I__937\ : Odrv4
    port map (
            O => \N__4329\,
            I => n1730
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__4326\,
            I => \N__4320\
        );

    \I__935\ : InMux
    port map (
            O => \N__4325\,
            I => \N__4314\
        );

    \I__934\ : InMux
    port map (
            O => \N__4324\,
            I => \N__4314\
        );

    \I__933\ : InMux
    port map (
            O => \N__4323\,
            I => \N__4311\
        );

    \I__932\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4306\
        );

    \I__931\ : InMux
    port map (
            O => \N__4319\,
            I => \N__4306\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4314\,
            I => i2c_cmd_cnt_1
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4311\,
            I => i2c_cmd_cnt_1
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4306\,
            I => i2c_cmd_cnt_1
        );

    \I__927\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4287\
        );

    \I__926\ : InMux
    port map (
            O => \N__4298\,
            I => \N__4287\
        );

    \I__925\ : InMux
    port map (
            O => \N__4297\,
            I => \N__4287\
        );

    \I__924\ : InMux
    port map (
            O => \N__4296\,
            I => \N__4280\
        );

    \I__923\ : InMux
    port map (
            O => \N__4295\,
            I => \N__4280\
        );

    \I__922\ : InMux
    port map (
            O => \N__4294\,
            I => \N__4280\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4287\,
            I => i2c_cmd_cnt_0
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4280\,
            I => i2c_cmd_cnt_0
        );

    \I__919\ : InMux
    port map (
            O => \N__4275\,
            I => \N__4271\
        );

    \I__918\ : InMux
    port map (
            O => \N__4274\,
            I => \N__4268\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4271\,
            I => \N__4265\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4268\,
            I => i2c_cmd_cnt_2
        );

    \I__915\ : Odrv4
    port map (
            O => \N__4265\,
            I => i2c_cmd_cnt_2
        );

    \I__914\ : ClkMux
    port map (
            O => \N__4260\,
            I => \N__4197\
        );

    \I__913\ : ClkMux
    port map (
            O => \N__4259\,
            I => \N__4197\
        );

    \I__912\ : ClkMux
    port map (
            O => \N__4258\,
            I => \N__4197\
        );

    \I__911\ : ClkMux
    port map (
            O => \N__4257\,
            I => \N__4197\
        );

    \I__910\ : ClkMux
    port map (
            O => \N__4256\,
            I => \N__4197\
        );

    \I__909\ : ClkMux
    port map (
            O => \N__4255\,
            I => \N__4197\
        );

    \I__908\ : ClkMux
    port map (
            O => \N__4254\,
            I => \N__4197\
        );

    \I__907\ : ClkMux
    port map (
            O => \N__4253\,
            I => \N__4197\
        );

    \I__906\ : ClkMux
    port map (
            O => \N__4252\,
            I => \N__4197\
        );

    \I__905\ : ClkMux
    port map (
            O => \N__4251\,
            I => \N__4197\
        );

    \I__904\ : ClkMux
    port map (
            O => \N__4250\,
            I => \N__4197\
        );

    \I__903\ : ClkMux
    port map (
            O => \N__4249\,
            I => \N__4197\
        );

    \I__902\ : ClkMux
    port map (
            O => \N__4248\,
            I => \N__4197\
        );

    \I__901\ : ClkMux
    port map (
            O => \N__4247\,
            I => \N__4197\
        );

    \I__900\ : ClkMux
    port map (
            O => \N__4246\,
            I => \N__4197\
        );

    \I__899\ : ClkMux
    port map (
            O => \N__4245\,
            I => \N__4197\
        );

    \I__898\ : ClkMux
    port map (
            O => \N__4244\,
            I => \N__4197\
        );

    \I__897\ : ClkMux
    port map (
            O => \N__4243\,
            I => \N__4197\
        );

    \I__896\ : ClkMux
    port map (
            O => \N__4242\,
            I => \N__4197\
        );

    \I__895\ : ClkMux
    port map (
            O => \N__4241\,
            I => \N__4197\
        );

    \I__894\ : ClkMux
    port map (
            O => \N__4240\,
            I => \N__4197\
        );

    \I__893\ : GlobalMux
    port map (
            O => \N__4197\,
            I => \N__4194\
        );

    \I__892\ : gio2CtrlBuf
    port map (
            O => \N__4194\,
            I => sysclk
        );

    \I__891\ : CEMux
    port map (
            O => \N__4191\,
            I => \N__4188\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4188\,
            I => \N__4185\
        );

    \I__889\ : Span4Mux_h
    port map (
            O => \N__4185\,
            I => \N__4182\
        );

    \I__888\ : Span4Mux_s3_h
    port map (
            O => \N__4182\,
            I => \N__4179\
        );

    \I__887\ : Odrv4
    port map (
            O => \N__4179\,
            I => n2956
        );

    \I__886\ : SRMux
    port map (
            O => \N__4176\,
            I => \N__4173\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4173\,
            I => \N__4170\
        );

    \I__884\ : Span4Mux_h
    port map (
            O => \N__4170\,
            I => \N__4167\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__4167\,
            I => n2016
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__4164\,
            I => \n25_cascade_\
        );

    \I__881\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4157\
        );

    \I__880\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4153\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4157\,
            I => \N__4150\
        );

    \I__878\ : InMux
    port map (
            O => \N__4156\,
            I => \N__4147\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4153\,
            I => \N__4142\
        );

    \I__876\ : Span4Mux_h
    port map (
            O => \N__4150\,
            I => \N__4142\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4147\,
            I => \N__4137\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__4142\,
            I => \N__4137\
        );

    \I__873\ : DummyBuf
    port map (
            O => \N__4137\,
            I => \hard0_SBDATo_2\
        );

    \I__872\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4131\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4131\,
            I => n2534
        );

    \I__870\ : InMux
    port map (
            O => \N__4128\,
            I => \N__4125\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4125\,
            I => \N__4122\
        );

    \I__868\ : Odrv4
    port map (
            O => \N__4122\,
            I => n4_adj_1
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__4119\,
            I => \n2840_cascade_\
        );

    \I__866\ : InMux
    port map (
            O => \N__4116\,
            I => \N__4113\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4113\,
            I => n2850
        );

    \I__864\ : CascadeMux
    port map (
            O => \N__4110\,
            I => \n29_cascade_\
        );

    \I__863\ : InMux
    port map (
            O => \N__4107\,
            I => \N__4104\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4104\,
            I => n26
        );

    \I__861\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4098\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4098\,
            I => n2958
        );

    \I__859\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4092\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4092\,
            I => \i2c_stat_7_N_205_2\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__4089\,
            I => \n2958_cascade_\
        );

    \I__856\ : InMux
    port map (
            O => \N__4086\,
            I => \N__4082\
        );

    \I__855\ : InMux
    port map (
            O => \N__4085\,
            I => \N__4079\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4082\,
            I => n20
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4079\,
            I => n20
        );

    \I__852\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4070\
        );

    \I__851\ : InMux
    port map (
            O => \N__4073\,
            I => \N__4067\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4070\,
            I => \N__4064\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4067\,
            I => cmd_decoded
        );

    \I__848\ : Odrv4
    port map (
            O => \N__4064\,
            I => cmd_decoded
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__4059\,
            I => \n2961_cascade_\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__4056\,
            I => \N__4053\
        );

    \I__845\ : InMux
    port map (
            O => \N__4053\,
            I => \N__4045\
        );

    \I__844\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4045\
        );

    \I__843\ : InMux
    port map (
            O => \N__4051\,
            I => \N__4042\
        );

    \I__842\ : InMux
    port map (
            O => \N__4050\,
            I => \N__4039\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4045\,
            I => \N__4036\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4042\,
            I => n2961
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4039\,
            I => n2961
        );

    \I__838\ : Odrv4
    port map (
            O => \N__4036\,
            I => n2961
        );

    \I__837\ : InMux
    port map (
            O => \N__4029\,
            I => \N__4026\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4026\,
            I => n2973
        );

    \I__835\ : InMux
    port map (
            O => \N__4023\,
            I => \N__4020\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4020\,
            I => n2962
        );

    \I__833\ : InMux
    port map (
            O => \N__4017\,
            I => \N__4014\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4014\,
            I => \N__4011\
        );

    \I__831\ : Span4Mux_s1_v
    port map (
            O => \N__4011\,
            I => \N__4006\
        );

    \I__830\ : InMux
    port map (
            O => \N__4010\,
            I => \N__4003\
        );

    \I__829\ : InMux
    port map (
            O => \N__4009\,
            I => \N__4000\
        );

    \I__828\ : Span4Mux_h
    port map (
            O => \N__4006\,
            I => \N__3997\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4003\,
            I => \N__3990\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4000\,
            I => \N__3990\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__3997\,
            I => \N__3990\
        );

    \I__824\ : DummyBuf
    port map (
            O => \N__3990\,
            I => \hard0_SBDATo_6\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__3987\,
            I => \i2c_stat_7_N_205_6_cascade_\
        );

    \I__822\ : InMux
    port map (
            O => \N__3984\,
            I => \N__3974\
        );

    \I__821\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3974\
        );

    \I__820\ : InMux
    port map (
            O => \N__3982\,
            I => \N__3974\
        );

    \I__819\ : InMux
    port map (
            O => \N__3981\,
            I => \N__3971\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__3974\,
            I => i2c_stat_6
        );

    \I__817\ : LocalMux
    port map (
            O => \N__3971\,
            I => i2c_stat_6
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__3966\,
            I => \N__3962\
        );

    \I__815\ : InMux
    port map (
            O => \N__3965\,
            I => \N__3957\
        );

    \I__814\ : InMux
    port map (
            O => \N__3962\,
            I => \N__3950\
        );

    \I__813\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3950\
        );

    \I__812\ : InMux
    port map (
            O => \N__3960\,
            I => \N__3950\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__3957\,
            I => i2c_cnt_1
        );

    \I__810\ : LocalMux
    port map (
            O => \N__3950\,
            I => i2c_cnt_1
        );

    \I__809\ : InMux
    port map (
            O => \N__3945\,
            I => \N__3939\
        );

    \I__808\ : InMux
    port map (
            O => \N__3944\,
            I => \N__3932\
        );

    \I__807\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3932\
        );

    \I__806\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3932\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__3939\,
            I => i2c_cnt_0
        );

    \I__804\ : LocalMux
    port map (
            O => \N__3932\,
            I => i2c_cnt_0
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__3927\,
            I => \n2534_cascade_\
        );

    \I__802\ : SRMux
    port map (
            O => \N__3924\,
            I => \N__3921\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__3921\,
            I => \N__3916\
        );

    \I__800\ : InMux
    port map (
            O => \N__3920\,
            I => \N__3911\
        );

    \I__799\ : InMux
    port map (
            O => \N__3919\,
            I => \N__3911\
        );

    \I__798\ : Span4Mux_v
    port map (
            O => \N__3916\,
            I => \N__3908\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__3911\,
            I => \N__3905\
        );

    \I__796\ : Odrv4
    port map (
            O => \N__3908\,
            I => n2959
        );

    \I__795\ : Odrv4
    port map (
            O => \N__3905\,
            I => n2959
        );

    \I__794\ : InMux
    port map (
            O => \N__3900\,
            I => \N__3897\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__3897\,
            I => n1887
        );

    \I__792\ : InMux
    port map (
            O => \N__3894\,
            I => \N__3888\
        );

    \I__791\ : InMux
    port map (
            O => \N__3893\,
            I => \N__3888\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__3888\,
            I => n4
        );

    \I__789\ : CEMux
    port map (
            O => \N__3885\,
            I => \N__3882\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__3882\,
            I => \N__3878\
        );

    \I__787\ : CEMux
    port map (
            O => \N__3881\,
            I => \N__3875\
        );

    \I__786\ : Span4Mux_s2_h
    port map (
            O => \N__3878\,
            I => \N__3870\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__3875\,
            I => \N__3870\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__3870\,
            I => n1779
        );

    \I__783\ : InMux
    port map (
            O => \N__3867\,
            I => \N__3861\
        );

    \I__782\ : InMux
    port map (
            O => \N__3866\,
            I => \N__3854\
        );

    \I__781\ : InMux
    port map (
            O => \N__3865\,
            I => \N__3854\
        );

    \I__780\ : InMux
    port map (
            O => \N__3864\,
            I => \N__3854\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__3861\,
            I => \N__3851\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__3854\,
            I => n2972
        );

    \I__777\ : Odrv4
    port map (
            O => \N__3851\,
            I => n2972
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__3846\,
            I => \n13_cascade_\
        );

    \I__775\ : CascadeMux
    port map (
            O => \N__3843\,
            I => \n4_adj_19_cascade_\
        );

    \I__774\ : DummyBuf
    port map (
            O => \N__3840\,
            I => \N__3837\
        );

    \I__773\ : InMux
    port map (
            O => \N__3837\,
            I => \N__3834\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__3834\,
            I => \N__3831\
        );

    \I__771\ : Span4Mux_s1_h
    port map (
            O => \N__3831\,
            I => \N__3827\
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__3830\,
            I => \N__3823\
        );

    \I__769\ : Span4Mux_h
    port map (
            O => \N__3827\,
            I => \N__3820\
        );

    \I__768\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3817\
        );

    \I__767\ : InMux
    port map (
            O => \N__3823\,
            I => \N__3814\
        );

    \I__766\ : Odrv4
    port map (
            O => \N__3820\,
            I => \hard_SBADRi_1\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__3817\,
            I => \hard_SBADRi_1\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__3814\,
            I => \hard_SBADRi_1\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__3807\,
            I => \n13_adj_4_cascade_\
        );

    \I__762\ : DummyBuf
    port map (
            O => \N__3804\,
            I => \N__3801\
        );

    \I__761\ : InMux
    port map (
            O => \N__3801\,
            I => \N__3798\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__3798\,
            I => \N__3795\
        );

    \I__759\ : Span4Mux_s1_h
    port map (
            O => \N__3795\,
            I => \N__3791\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__3794\,
            I => \N__3787\
        );

    \I__757\ : Span4Mux_h
    port map (
            O => \N__3791\,
            I => \N__3784\
        );

    \I__756\ : InMux
    port map (
            O => \N__3790\,
            I => \N__3781\
        );

    \I__755\ : InMux
    port map (
            O => \N__3787\,
            I => \N__3778\
        );

    \I__754\ : Odrv4
    port map (
            O => \N__3784\,
            I => \hard_SBDATi_7\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__3781\,
            I => \hard_SBDATi_7\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__3778\,
            I => \hard_SBDATi_7\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__3771\,
            I => \n2974_cascade_\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__3768\,
            I => \n2970_cascade_\
        );

    \I__749\ : DummyBuf
    port map (
            O => \N__3765\,
            I => \N__3762\
        );

    \I__748\ : InMux
    port map (
            O => \N__3762\,
            I => \N__3758\
        );

    \I__747\ : InMux
    port map (
            O => \N__3761\,
            I => \N__3755\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__3758\,
            I => \N__3752\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3755\,
            I => \hard_SBSTBi\
        );

    \I__744\ : Odrv12
    port map (
            O => \N__3752\,
            I => \hard_SBSTBi\
        );

    \I__743\ : InMux
    port map (
            O => \N__3747\,
            I => \N__3744\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__3744\,
            I => n31
        );

    \I__741\ : InMux
    port map (
            O => \N__3741\,
            I => \N__3738\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3738\,
            I => n2970
        );

    \I__739\ : InMux
    port map (
            O => \N__3735\,
            I => \N__3731\
        );

    \I__738\ : InMux
    port map (
            O => \N__3734\,
            I => \N__3728\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3731\,
            I => \N__3725\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3728\,
            I => n2243
        );

    \I__735\ : Odrv4
    port map (
            O => \N__3725\,
            I => n2243
        );

    \I__734\ : CascadeMux
    port map (
            O => \N__3720\,
            I => \n17_cascade_\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__3717\,
            I => \n1887_cascade_\
        );

    \I__732\ : InMux
    port map (
            O => \N__3714\,
            I => \N__3711\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__3711\,
            I => n1852
        );

    \I__730\ : InMux
    port map (
            O => \N__3708\,
            I => \N__3705\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3705\,
            I => n22_adj_9
        );

    \I__728\ : InMux
    port map (
            O => \N__3702\,
            I => \N__3698\
        );

    \I__727\ : InMux
    port map (
            O => \N__3701\,
            I => \N__3695\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__3698\,
            I => n2971
        );

    \I__725\ : LocalMux
    port map (
            O => \N__3695\,
            I => n2971
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__3690\,
            I => \n13_adj_6_cascade_\
        );

    \I__723\ : DummyBuf
    port map (
            O => \N__3687\,
            I => \N__3684\
        );

    \I__722\ : InMux
    port map (
            O => \N__3684\,
            I => \N__3681\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__3681\,
            I => \N__3677\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__3680\,
            I => \N__3673\
        );

    \I__719\ : Span4Mux_h
    port map (
            O => \N__3677\,
            I => \N__3670\
        );

    \I__718\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3665\
        );

    \I__717\ : InMux
    port map (
            O => \N__3673\,
            I => \N__3665\
        );

    \I__716\ : Odrv4
    port map (
            O => \N__3670\,
            I => \hard_SBDATi_4\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3665\,
            I => \hard_SBDATi_4\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__3660\,
            I => \n12_cascade_\
        );

    \I__713\ : DummyBuf
    port map (
            O => \N__3657\,
            I => \N__3654\
        );

    \I__712\ : InMux
    port map (
            O => \N__3654\,
            I => \N__3651\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3651\,
            I => \N__3647\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__3650\,
            I => \N__3643\
        );

    \I__709\ : Span4Mux_s1_v
    port map (
            O => \N__3647\,
            I => \N__3640\
        );

    \I__708\ : InMux
    port map (
            O => \N__3646\,
            I => \N__3635\
        );

    \I__707\ : InMux
    port map (
            O => \N__3643\,
            I => \N__3635\
        );

    \I__706\ : Odrv4
    port map (
            O => \N__3640\,
            I => \hard_SBDATi_2\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3635\,
            I => \hard_SBDATi_2\
        );

    \I__704\ : InMux
    port map (
            O => \N__3630\,
            I => \N__3627\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3627\,
            I => n15
        );

    \I__702\ : CascadeMux
    port map (
            O => \N__3624\,
            I => \n2824_cascade_\
        );

    \I__701\ : DummyBuf
    port map (
            O => \N__3621\,
            I => \N__3618\
        );

    \I__700\ : InMux
    port map (
            O => \N__3618\,
            I => \N__3615\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3615\,
            I => \N__3611\
        );

    \I__698\ : InMux
    port map (
            O => \N__3614\,
            I => \N__3608\
        );

    \I__697\ : Span12Mux_s4_h
    port map (
            O => \N__3611\,
            I => \N__3605\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3608\,
            I => \hard_SBADRi_3\
        );

    \I__695\ : Odrv12
    port map (
            O => \N__3605\,
            I => \hard_SBADRi_3\
        );

    \I__694\ : InMux
    port map (
            O => \N__3600\,
            I => \N__3597\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3597\,
            I => \N__3593\
        );

    \I__692\ : DummyBuf
    port map (
            O => \N__3596\,
            I => \N__3590\
        );

    \I__691\ : Glb2LocalMux
    port map (
            O => \N__3593\,
            I => \N__3585\
        );

    \I__690\ : ClkMux
    port map (
            O => \N__3590\,
            I => \N__3585\
        );

    \I__689\ : GlobalMux
    port map (
            O => \N__3585\,
            I => \N__3582\
        );

    \I__688\ : DummyBuf
    port map (
            O => \N__3582\,
            I => n2981
        );

    \I__687\ : IoInMux
    port map (
            O => \N__3579\,
            I => \N__3576\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3576\,
            I => \N__3573\
        );

    \I__685\ : IoSpan4Mux
    port map (
            O => \N__3573\,
            I => \N__3570\
        );

    \I__684\ : Odrv4
    port map (
            O => \N__3570\,
            I => \GB_BUFFER_n2981_THRU_CO\
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__3567\,
            I => \n2960_cascade_\
        );

    \I__682\ : DummyBuf
    port map (
            O => \N__3564\,
            I => \N__3561\
        );

    \I__681\ : InMux
    port map (
            O => \N__3561\,
            I => \N__3557\
        );

    \I__680\ : InMux
    port map (
            O => \N__3560\,
            I => \N__3554\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3557\,
            I => \N__3551\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3554\,
            I => \hard_SBWRi\
        );

    \I__677\ : Odrv12
    port map (
            O => \N__3551\,
            I => \hard_SBWRi\
        );

    \I__676\ : DummyBuf
    port map (
            O => \N__3546\,
            I => \N__3542\
        );

    \I__675\ : CascadeMux
    port map (
            O => \N__3545\,
            I => \N__3539\
        );

    \I__674\ : InMux
    port map (
            O => \N__3542\,
            I => \N__3536\
        );

    \I__673\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3533\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3536\,
            I => \N__3530\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3533\,
            I => \hard_SBADRi_0\
        );

    \I__670\ : Odrv12
    port map (
            O => \N__3530\,
            I => \hard_SBADRi_0\
        );

    \I__669\ : CascadeMux
    port map (
            O => \N__3525\,
            I => \n12_adj_7_cascade_\
        );

    \I__668\ : DummyBuf
    port map (
            O => \N__3522\,
            I => \N__3519\
        );

    \I__667\ : InMux
    port map (
            O => \N__3519\,
            I => \N__3515\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__3518\,
            I => \N__3511\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3515\,
            I => \N__3508\
        );

    \I__664\ : InMux
    port map (
            O => \N__3514\,
            I => \N__3503\
        );

    \I__663\ : InMux
    port map (
            O => \N__3511\,
            I => \N__3503\
        );

    \I__662\ : Odrv12
    port map (
            O => \N__3508\,
            I => \hard_SBADRi_2\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3503\,
            I => \hard_SBADRi_2\
        );

    \I__660\ : InMux
    port map (
            O => \N__3498\,
            I => \N__3495\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3495\,
            I => n8_adj_10
        );

    \I__658\ : InMux
    port map (
            O => \N__3492\,
            I => \N__3489\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3489\,
            I => \N__3485\
        );

    \I__656\ : InMux
    port map (
            O => \N__3488\,
            I => \N__3482\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__3485\,
            I => n2881
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3482\,
            I => n2881
        );

    \I__653\ : InMux
    port map (
            O => \N__3477\,
            I => \N__3474\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3474\,
            I => n14_adj_14
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__3471\,
            I => \n104_cascade_\
        );

    \I__650\ : InMux
    port map (
            O => \N__3468\,
            I => \N__3465\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3465\,
            I => \N__3457\
        );

    \I__648\ : InMux
    port map (
            O => \N__3464\,
            I => \N__3450\
        );

    \I__647\ : InMux
    port map (
            O => \N__3463\,
            I => \N__3450\
        );

    \I__646\ : InMux
    port map (
            O => \N__3462\,
            I => \N__3450\
        );

    \I__645\ : InMux
    port map (
            O => \N__3461\,
            I => \N__3445\
        );

    \I__644\ : InMux
    port map (
            O => \N__3460\,
            I => \N__3445\
        );

    \I__643\ : Span4Mux_v
    port map (
            O => \N__3457\,
            I => \N__3442\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3450\,
            I => n105
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3445\,
            I => n105
        );

    \I__640\ : Odrv4
    port map (
            O => \N__3442\,
            I => n105
        );

    \I__639\ : SRMux
    port map (
            O => \N__3435\,
            I => \N__3432\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3432\,
            I => \N__3429\
        );

    \I__637\ : Odrv4
    port map (
            O => \N__3429\,
            I => n1921
        );

    \I__636\ : InMux
    port map (
            O => \N__3426\,
            I => \N__3423\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3423\,
            I => \N__3418\
        );

    \I__634\ : InMux
    port map (
            O => \N__3422\,
            I => \N__3413\
        );

    \I__633\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3413\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__3418\,
            I => \PWM_duty_7\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3413\,
            I => \PWM_duty_7\
        );

    \I__630\ : InMux
    port map (
            O => \N__3408\,
            I => \N__3402\
        );

    \I__629\ : InMux
    port map (
            O => \N__3407\,
            I => \N__3399\
        );

    \I__628\ : InMux
    port map (
            O => \N__3406\,
            I => \N__3396\
        );

    \I__627\ : InMux
    port map (
            O => \N__3405\,
            I => \N__3393\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3402\,
            I => \PWM_cnt_7\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3399\,
            I => \PWM_cnt_7\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3396\,
            I => \PWM_cnt_7\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3393\,
            I => \PWM_cnt_7\
        );

    \I__622\ : InMux
    port map (
            O => \N__3384\,
            I => \N__3380\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__3383\,
            I => \N__3377\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3380\,
            I => \N__3374\
        );

    \I__619\ : InMux
    port map (
            O => \N__3377\,
            I => \N__3371\
        );

    \I__618\ : Odrv12
    port map (
            O => \N__3374\,
            I => n2969
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3371\,
            I => n2969
        );

    \I__616\ : InMux
    port map (
            O => \N__3366\,
            I => \N__3361\
        );

    \I__615\ : InMux
    port map (
            O => \N__3365\,
            I => \N__3358\
        );

    \I__614\ : InMux
    port map (
            O => \N__3364\,
            I => \N__3355\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3361\,
            I => drv_clk_counter_4
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3358\,
            I => drv_clk_counter_4
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3355\,
            I => drv_clk_counter_4
        );

    \I__610\ : InMux
    port map (
            O => \N__3348\,
            I => \N__3343\
        );

    \I__609\ : InMux
    port map (
            O => \N__3347\,
            I => \N__3340\
        );

    \I__608\ : InMux
    port map (
            O => \N__3346\,
            I => \N__3337\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3343\,
            I => drv_clk_counter_1
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3340\,
            I => drv_clk_counter_1
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3337\,
            I => drv_clk_counter_1
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__3330\,
            I => \N__3326\
        );

    \I__603\ : InMux
    port map (
            O => \N__3329\,
            I => \N__3323\
        );

    \I__602\ : InMux
    port map (
            O => \N__3326\,
            I => \N__3320\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3323\,
            I => drv_clk_counter_0
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3320\,
            I => drv_clk_counter_0
        );

    \I__599\ : InMux
    port map (
            O => \N__3315\,
            I => \N__3310\
        );

    \I__598\ : InMux
    port map (
            O => \N__3314\,
            I => \N__3307\
        );

    \I__597\ : InMux
    port map (
            O => \N__3313\,
            I => \N__3304\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3310\,
            I => drv_clk_counter_8
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3307\,
            I => drv_clk_counter_8
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3304\,
            I => drv_clk_counter_8
        );

    \I__593\ : InMux
    port map (
            O => \N__3297\,
            I => \N__3292\
        );

    \I__592\ : InMux
    port map (
            O => \N__3296\,
            I => \N__3289\
        );

    \I__591\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3286\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3292\,
            I => drv_clk_counter_5
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3289\,
            I => drv_clk_counter_5
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3286\,
            I => drv_clk_counter_5
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__3279\,
            I => \n2810_cascade_\
        );

    \I__586\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3273\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3273\,
            I => \N__3269\
        );

    \I__584\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3266\
        );

    \I__583\ : Odrv4
    port map (
            O => \N__3269\,
            I => n2819
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3266\,
            I => n2819
        );

    \I__581\ : InMux
    port map (
            O => \N__3261\,
            I => \N__3250\
        );

    \I__580\ : InMux
    port map (
            O => \N__3260\,
            I => \N__3250\
        );

    \I__579\ : InMux
    port map (
            O => \N__3259\,
            I => \N__3250\
        );

    \I__578\ : InMux
    port map (
            O => \N__3258\,
            I => \N__3244\
        );

    \I__577\ : InMux
    port map (
            O => \N__3257\,
            I => \N__3244\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3250\,
            I => \N__3239\
        );

    \I__575\ : InMux
    port map (
            O => \N__3249\,
            I => \N__3236\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__3244\,
            I => \N__3233\
        );

    \I__573\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3230\
        );

    \I__572\ : InMux
    port map (
            O => \N__3242\,
            I => \N__3227\
        );

    \I__571\ : Span4Mux_s2_h
    port map (
            O => \N__3239\,
            I => \N__3224\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3236\,
            I => \N__3219\
        );

    \I__569\ : Span4Mux_s3_h
    port map (
            O => \N__3233\,
            I => \N__3219\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3230\,
            I => motor_on
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3227\,
            I => motor_on
        );

    \I__566\ : Odrv4
    port map (
            O => \N__3224\,
            I => motor_on
        );

    \I__565\ : Odrv4
    port map (
            O => \N__3219\,
            I => motor_on
        );

    \I__564\ : InMux
    port map (
            O => \N__3210\,
            I => \N__3205\
        );

    \I__563\ : InMux
    port map (
            O => \N__3209\,
            I => \N__3202\
        );

    \I__562\ : InMux
    port map (
            O => \N__3208\,
            I => \N__3199\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3205\,
            I => \N__3196\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3202\,
            I => drv_clk_counter_10
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3199\,
            I => drv_clk_counter_10
        );

    \I__558\ : Odrv4
    port map (
            O => \N__3196\,
            I => drv_clk_counter_10
        );

    \I__557\ : CascadeMux
    port map (
            O => \N__3189\,
            I => \n2820_cascade_\
        );

    \I__556\ : InMux
    port map (
            O => \N__3186\,
            I => \N__3181\
        );

    \I__555\ : InMux
    port map (
            O => \N__3185\,
            I => \N__3178\
        );

    \I__554\ : InMux
    port map (
            O => \N__3184\,
            I => \N__3175\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3181\,
            I => drv_clk_counter_9
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3178\,
            I => drv_clk_counter_9
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3175\,
            I => drv_clk_counter_9
        );

    \I__550\ : SRMux
    port map (
            O => \N__3168\,
            I => \N__3165\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3165\,
            I => \N__3161\
        );

    \I__548\ : SRMux
    port map (
            O => \N__3164\,
            I => \N__3158\
        );

    \I__547\ : Span4Mux_s2_h
    port map (
            O => \N__3161\,
            I => \N__3155\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3158\,
            I => \N__3152\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__3155\,
            I => n953
        );

    \I__544\ : Odrv4
    port map (
            O => \N__3152\,
            I => n953
        );

    \I__543\ : InMux
    port map (
            O => \N__3147\,
            I => \N__3142\
        );

    \I__542\ : InMux
    port map (
            O => \N__3146\,
            I => \N__3139\
        );

    \I__541\ : InMux
    port map (
            O => \N__3145\,
            I => \N__3136\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__3142\,
            I => drv_clk_counter_2
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3139\,
            I => drv_clk_counter_2
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3136\,
            I => drv_clk_counter_2
        );

    \I__537\ : InMux
    port map (
            O => \N__3129\,
            I => \N__3124\
        );

    \I__536\ : InMux
    port map (
            O => \N__3128\,
            I => \N__3121\
        );

    \I__535\ : InMux
    port map (
            O => \N__3127\,
            I => \N__3118\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3124\,
            I => drv_clk_counter_3
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3121\,
            I => drv_clk_counter_3
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3118\,
            I => drv_clk_counter_3
        );

    \I__531\ : InMux
    port map (
            O => \N__3111\,
            I => \N__3108\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3108\,
            I => n2963
        );

    \I__529\ : InMux
    port map (
            O => \N__3105\,
            I => \N__3099\
        );

    \I__528\ : InMux
    port map (
            O => \N__3104\,
            I => \N__3099\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3099\,
            I => n2247
        );

    \I__526\ : CascadeMux
    port map (
            O => \N__3096\,
            I => \n2250_cascade_\
        );

    \I__525\ : InMux
    port map (
            O => \N__3093\,
            I => \N__3086\
        );

    \I__524\ : InMux
    port map (
            O => \N__3092\,
            I => \N__3086\
        );

    \I__523\ : InMux
    port map (
            O => \N__3091\,
            I => \N__3083\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3086\,
            I => i2c_cmd_0_1
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3083\,
            I => i2c_cmd_0_1
        );

    \I__520\ : InMux
    port map (
            O => \N__3078\,
            I => \N__3069\
        );

    \I__519\ : InMux
    port map (
            O => \N__3077\,
            I => \N__3069\
        );

    \I__518\ : InMux
    port map (
            O => \N__3076\,
            I => \N__3069\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3069\,
            I => \N__3066\
        );

    \I__516\ : Odrv4
    port map (
            O => \N__3066\,
            I => i2c_cmd_0_4
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__3063\,
            I => \N__3059\
        );

    \I__514\ : InMux
    port map (
            O => \N__3062\,
            I => \N__3051\
        );

    \I__513\ : InMux
    port map (
            O => \N__3059\,
            I => \N__3051\
        );

    \I__512\ : InMux
    port map (
            O => \N__3058\,
            I => \N__3051\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3051\,
            I => i2c_cmd_0_0
        );

    \I__510\ : InMux
    port map (
            O => \N__3048\,
            I => \N__3045\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3045\,
            I => n2858
        );

    \I__508\ : CEMux
    port map (
            O => \N__3042\,
            I => \N__3039\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3039\,
            I => \N__3036\
        );

    \I__506\ : Odrv4
    port map (
            O => \N__3036\,
            I => n1778
        );

    \I__505\ : InMux
    port map (
            O => \N__3033\,
            I => \N__3028\
        );

    \I__504\ : InMux
    port map (
            O => \N__3032\,
            I => \N__3025\
        );

    \I__503\ : InMux
    port map (
            O => \N__3031\,
            I => \N__3022\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3028\,
            I => \PWM_duty_5\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3025\,
            I => \PWM_duty_5\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3022\,
            I => \PWM_duty_5\
        );

    \I__499\ : InMux
    port map (
            O => \N__3015\,
            I => \N__3011\
        );

    \I__498\ : InMux
    port map (
            O => \N__3014\,
            I => \N__3008\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3011\,
            I => n2968
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3008\,
            I => n2968
        );

    \I__495\ : InMux
    port map (
            O => \N__3003\,
            I => \N__3000\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3000\,
            I => n2883
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__2997\,
            I => \n2883_cascade_\
        );

    \I__492\ : InMux
    port map (
            O => \N__2994\,
            I => \N__2990\
        );

    \I__491\ : InMux
    port map (
            O => \N__2993\,
            I => \N__2987\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__2990\,
            I => \PWM_duty_0\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__2987\,
            I => \PWM_duty_0\
        );

    \I__488\ : InMux
    port map (
            O => \N__2982\,
            I => \N__2977\
        );

    \I__487\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2974\
        );

    \I__486\ : InMux
    port map (
            O => \N__2980\,
            I => \N__2971\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__2977\,
            I => \PWM_cnt_1\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__2974\,
            I => \PWM_cnt_1\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__2971\,
            I => \PWM_cnt_1\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__2964\,
            I => \N__2959\
        );

    \I__481\ : CascadeMux
    port map (
            O => \N__2963\,
            I => \N__2956\
        );

    \I__480\ : InMux
    port map (
            O => \N__2962\,
            I => \N__2953\
        );

    \I__479\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2950\
        );

    \I__478\ : InMux
    port map (
            O => \N__2956\,
            I => \N__2947\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__2953\,
            I => \PWM_cnt_0\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__2950\,
            I => \PWM_cnt_0\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__2947\,
            I => \PWM_cnt_0\
        );

    \I__474\ : InMux
    port map (
            O => \N__2940\,
            I => \N__2936\
        );

    \I__473\ : InMux
    port map (
            O => \N__2939\,
            I => \N__2933\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__2936\,
            I => \PWM_duty_1\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__2933\,
            I => \PWM_duty_1\
        );

    \I__470\ : InMux
    port map (
            O => \N__2928\,
            I => \N__2925\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2925\,
            I => n4_adj_17
        );

    \I__468\ : InMux
    port map (
            O => \N__2922\,
            I => \N__2917\
        );

    \I__467\ : InMux
    port map (
            O => \N__2921\,
            I => \N__2914\
        );

    \I__466\ : InMux
    port map (
            O => \N__2920\,
            I => \N__2911\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__2917\,
            I => \N__2908\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2914\,
            I => \PWM_duty_6\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2911\,
            I => \PWM_duty_6\
        );

    \I__462\ : Odrv4
    port map (
            O => \N__2908\,
            I => \PWM_duty_6\
        );

    \I__461\ : InMux
    port map (
            O => \N__2901\,
            I => \N__2895\
        );

    \I__460\ : InMux
    port map (
            O => \N__2900\,
            I => \N__2892\
        );

    \I__459\ : InMux
    port map (
            O => \N__2899\,
            I => \N__2889\
        );

    \I__458\ : InMux
    port map (
            O => \N__2898\,
            I => \N__2886\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__2895\,
            I => \PWM_cnt_6\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__2892\,
            I => \PWM_cnt_6\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__2889\,
            I => \PWM_cnt_6\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2886\,
            I => \PWM_cnt_6\
        );

    \I__453\ : InMux
    port map (
            O => \N__2877\,
            I => \N__2871\
        );

    \I__452\ : InMux
    port map (
            O => \N__2876\,
            I => \N__2868\
        );

    \I__451\ : InMux
    port map (
            O => \N__2875\,
            I => \N__2863\
        );

    \I__450\ : InMux
    port map (
            O => \N__2874\,
            I => \N__2863\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2871\,
            I => \PWM_cnt_5\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2868\,
            I => \PWM_cnt_5\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2863\,
            I => \PWM_cnt_5\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__2856\,
            I => \n10_cascade_\
        );

    \I__445\ : InMux
    port map (
            O => \N__2853\,
            I => \N__2850\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2850\,
            I => n12_adj_13
        );

    \I__443\ : CascadeMux
    port map (
            O => \N__2847\,
            I => \n2838_cascade_\
        );

    \I__442\ : InMux
    port map (
            O => \N__2844\,
            I => \N__2838\
        );

    \I__441\ : InMux
    port map (
            O => \N__2843\,
            I => \N__2838\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2838\,
            I => i2c_cmd_0_5
        );

    \I__439\ : InMux
    port map (
            O => \N__2835\,
            I => \N__2831\
        );

    \I__438\ : InMux
    port map (
            O => \N__2834\,
            I => \N__2828\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2831\,
            I => i2c_cmd_0_6
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2828\,
            I => i2c_cmd_0_6
        );

    \I__435\ : InMux
    port map (
            O => \N__2823\,
            I => \N__2817\
        );

    \I__434\ : InMux
    port map (
            O => \N__2822\,
            I => \N__2817\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__2817\,
            I => i2c_cmd_0_3
        );

    \I__432\ : CascadeMux
    port map (
            O => \N__2814\,
            I => \n6_adj_8_cascade_\
        );

    \I__431\ : InMux
    port map (
            O => \N__2811\,
            I => \N__2805\
        );

    \I__430\ : InMux
    port map (
            O => \N__2810\,
            I => \N__2805\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2805\,
            I => i2c_cmd_0_7
        );

    \I__428\ : InMux
    port map (
            O => \N__2802\,
            I => \N__2796\
        );

    \I__427\ : InMux
    port map (
            O => \N__2801\,
            I => \N__2796\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2796\,
            I => i2c_cmd_0_2
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__2793\,
            I => \N__2790\
        );

    \I__424\ : InMux
    port map (
            O => \N__2790\,
            I => \N__2787\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2787\,
            I => \N__2784\
        );

    \I__422\ : Odrv4
    port map (
            O => \N__2784\,
            I => n10_adj_2
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__2781\,
            I => \n17_adj_18_cascade_\
        );

    \I__420\ : InMux
    port map (
            O => \N__2778\,
            I => \N__2773\
        );

    \I__419\ : InMux
    port map (
            O => \N__2777\,
            I => \N__2770\
        );

    \I__418\ : InMux
    port map (
            O => \N__2776\,
            I => \N__2767\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2773\,
            I => \PWM_cnt_2\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2770\,
            I => \PWM_cnt_2\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2767\,
            I => \PWM_cnt_2\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__2760\,
            I => \N__2755\
        );

    \I__413\ : InMux
    port map (
            O => \N__2759\,
            I => \N__2751\
        );

    \I__412\ : InMux
    port map (
            O => \N__2758\,
            I => \N__2748\
        );

    \I__411\ : InMux
    port map (
            O => \N__2755\,
            I => \N__2743\
        );

    \I__410\ : InMux
    port map (
            O => \N__2754\,
            I => \N__2743\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2751\,
            I => \PWM_cnt_3\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2748\,
            I => \PWM_cnt_3\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2743\,
            I => \PWM_cnt_3\
        );

    \I__406\ : InMux
    port map (
            O => \N__2736\,
            I => \N__2731\
        );

    \I__405\ : InMux
    port map (
            O => \N__2735\,
            I => \N__2726\
        );

    \I__404\ : InMux
    port map (
            O => \N__2734\,
            I => \N__2726\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2731\,
            I => \PWM_duty_3\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2726\,
            I => \PWM_duty_3\
        );

    \I__401\ : InMux
    port map (
            O => \N__2721\,
            I => \N__2716\
        );

    \I__400\ : InMux
    port map (
            O => \N__2720\,
            I => \N__2711\
        );

    \I__399\ : InMux
    port map (
            O => \N__2719\,
            I => \N__2711\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2716\,
            I => \PWM_duty_4\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2711\,
            I => \PWM_duty_4\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__2706\,
            I => \n6_adj_5_cascade_\
        );

    \I__395\ : InMux
    port map (
            O => \N__2703\,
            I => \N__2697\
        );

    \I__394\ : InMux
    port map (
            O => \N__2702\,
            I => \N__2694\
        );

    \I__393\ : InMux
    port map (
            O => \N__2701\,
            I => \N__2689\
        );

    \I__392\ : InMux
    port map (
            O => \N__2700\,
            I => \N__2689\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2697\,
            I => \PWM_cnt_4\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__2694\,
            I => \PWM_cnt_4\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2689\,
            I => \PWM_cnt_4\
        );

    \I__388\ : InMux
    port map (
            O => \N__2682\,
            I => n2523
        );

    \I__387\ : InMux
    port map (
            O => \N__2679\,
            I => n2524
        );

    \I__386\ : InMux
    port map (
            O => \N__2676\,
            I => n2525
        );

    \I__385\ : InMux
    port map (
            O => \N__2673\,
            I => \N__2669\
        );

    \I__384\ : InMux
    port map (
            O => \N__2672\,
            I => \N__2666\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2669\,
            I => drv_clk_counter_6
        );

    \I__382\ : LocalMux
    port map (
            O => \N__2666\,
            I => drv_clk_counter_6
        );

    \I__381\ : InMux
    port map (
            O => \N__2661\,
            I => n2526
        );

    \I__380\ : InMux
    port map (
            O => \N__2658\,
            I => \N__2654\
        );

    \I__379\ : InMux
    port map (
            O => \N__2657\,
            I => \N__2651\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2654\,
            I => drv_clk_counter_7
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2651\,
            I => drv_clk_counter_7
        );

    \I__376\ : InMux
    port map (
            O => \N__2646\,
            I => n2527
        );

    \I__375\ : InMux
    port map (
            O => \N__2643\,
            I => \bfn_1_7_0_\
        );

    \I__374\ : InMux
    port map (
            O => \N__2640\,
            I => n2529
        );

    \I__373\ : InMux
    port map (
            O => \N__2637\,
            I => n2530
        );

    \I__372\ : CascadeMux
    port map (
            O => \N__2634\,
            I => \n12_adj_11_cascade_\
        );

    \I__371\ : InMux
    port map (
            O => \N__2631\,
            I => \N__2628\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2628\,
            I => n4_adj_15
        );

    \I__369\ : InMux
    port map (
            O => \N__2625\,
            I => \N__2622\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2622\,
            I => n8
        );

    \I__367\ : CascadeMux
    port map (
            O => \N__2619\,
            I => \n14_cascade_\
        );

    \I__366\ : CascadeMux
    port map (
            O => \N__2616\,
            I => \N__2612\
        );

    \I__365\ : InMux
    port map (
            O => \N__2615\,
            I => \N__2608\
        );

    \I__364\ : InMux
    port map (
            O => \N__2612\,
            I => \N__2603\
        );

    \I__363\ : InMux
    port map (
            O => \N__2611\,
            I => \N__2603\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2608\,
            I => n2012
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2603\,
            I => n2012
        );

    \I__360\ : CEMux
    port map (
            O => \N__2598\,
            I => \N__2595\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2595\,
            I => \N__2592\
        );

    \I__358\ : Odrv12
    port map (
            O => \N__2592\,
            I => n2955
        );

    \I__357\ : CascadeMux
    port map (
            O => \N__2589\,
            I => \N__2585\
        );

    \I__356\ : InMux
    port map (
            O => \N__2588\,
            I => \N__2581\
        );

    \I__355\ : InMux
    port map (
            O => \N__2585\,
            I => \N__2575\
        );

    \I__354\ : InMux
    port map (
            O => \N__2584\,
            I => \N__2575\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2581\,
            I => \N__2571\
        );

    \I__352\ : InMux
    port map (
            O => \N__2580\,
            I => \N__2568\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2575\,
            I => \N__2565\
        );

    \I__350\ : InMux
    port map (
            O => \N__2574\,
            I => \N__2562\
        );

    \I__349\ : Odrv4
    port map (
            O => \N__2571\,
            I => drv_cnt_1
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2568\,
            I => drv_cnt_1
        );

    \I__347\ : Odrv4
    port map (
            O => \N__2565\,
            I => drv_cnt_1
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2562\,
            I => drv_cnt_1
        );

    \I__345\ : InMux
    port map (
            O => \N__2553\,
            I => \N__2546\
        );

    \I__344\ : InMux
    port map (
            O => \N__2552\,
            I => \N__2546\
        );

    \I__343\ : InMux
    port map (
            O => \N__2551\,
            I => \N__2540\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2546\,
            I => \N__2537\
        );

    \I__341\ : InMux
    port map (
            O => \N__2545\,
            I => \N__2532\
        );

    \I__340\ : InMux
    port map (
            O => \N__2544\,
            I => \N__2532\
        );

    \I__339\ : InMux
    port map (
            O => \N__2543\,
            I => \N__2529\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2540\,
            I => drv_cnt_0
        );

    \I__337\ : Odrv4
    port map (
            O => \N__2537\,
            I => drv_cnt_0
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2532\,
            I => drv_cnt_0
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2529\,
            I => drv_cnt_0
        );

    \I__334\ : CascadeMux
    port map (
            O => \N__2520\,
            I => \n2955_cascade_\
        );

    \I__333\ : InMux
    port map (
            O => \N__2517\,
            I => \N__2509\
        );

    \I__332\ : InMux
    port map (
            O => \N__2516\,
            I => \N__2509\
        );

    \I__331\ : InMux
    port map (
            O => \N__2515\,
            I => \N__2505\
        );

    \I__330\ : InMux
    port map (
            O => \N__2514\,
            I => \N__2502\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2509\,
            I => \N__2499\
        );

    \I__328\ : InMux
    port map (
            O => \N__2508\,
            I => \N__2496\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2505\,
            I => drv_cnt_2
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2502\,
            I => drv_cnt_2
        );

    \I__325\ : Odrv4
    port map (
            O => \N__2499\,
            I => drv_cnt_2
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2496\,
            I => drv_cnt_2
        );

    \I__323\ : InMux
    port map (
            O => \N__2487\,
            I => \bfn_1_6_0_\
        );

    \I__322\ : InMux
    port map (
            O => \N__2484\,
            I => n2521
        );

    \I__321\ : InMux
    port map (
            O => \N__2481\,
            I => n2522
        );

    \I__320\ : InMux
    port map (
            O => \N__2478\,
            I => n2514
        );

    \I__319\ : InMux
    port map (
            O => \N__2475\,
            I => n2515
        );

    \I__318\ : InMux
    port map (
            O => \N__2472\,
            I => n2516
        );

    \I__317\ : InMux
    port map (
            O => \N__2469\,
            I => n2517
        );

    \I__316\ : InMux
    port map (
            O => \N__2466\,
            I => n2518
        );

    \I__315\ : InMux
    port map (
            O => \N__2463\,
            I => n2519
        );

    \I__314\ : InMux
    port map (
            O => \N__2460\,
            I => n2520
        );

    \I__313\ : CEMux
    port map (
            O => \N__2457\,
            I => \N__2454\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2454\,
            I => \N__2451\
        );

    \I__311\ : Odrv12
    port map (
            O => \N__2451\,
            I => n1831
        );

    \I__310\ : InMux
    port map (
            O => \N__2448\,
            I => \N__2445\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2445\,
            I => \N__2442\
        );

    \I__308\ : Odrv4
    port map (
            O => \N__2442\,
            I => i2c_cmd_1_0
        );

    \I__307\ : InMux
    port map (
            O => \N__2439\,
            I => \N__2436\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2436\,
            I => \N__2433\
        );

    \I__305\ : Odrv4
    port map (
            O => \N__2433\,
            I => i2c_cmd_1_1
        );

    \I__304\ : InMux
    port map (
            O => \N__2430\,
            I => \N__2427\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2427\,
            I => \N__2424\
        );

    \I__302\ : Odrv4
    port map (
            O => \N__2424\,
            I => i2c_cmd_1_2
        );

    \I__301\ : InMux
    port map (
            O => \N__2421\,
            I => \N__2415\
        );

    \I__300\ : InMux
    port map (
            O => \N__2420\,
            I => \N__2415\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2415\,
            I => \PWM_duty_2\
        );

    \I__298\ : InMux
    port map (
            O => \N__2412\,
            I => \N__2409\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2409\,
            I => \N__2406\
        );

    \I__296\ : Odrv4
    port map (
            O => \N__2406\,
            I => i2c_cmd_1_5
        );

    \I__295\ : InMux
    port map (
            O => \N__2403\,
            I => \N__2400\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2400\,
            I => \N__2397\
        );

    \I__293\ : Odrv4
    port map (
            O => \N__2397\,
            I => i2c_cmd_1_6
        );

    \I__292\ : InMux
    port map (
            O => \N__2394\,
            I => \N__2391\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2391\,
            I => \N__2388\
        );

    \I__290\ : Odrv4
    port map (
            O => \N__2388\,
            I => i2c_cmd_1_7
        );

    \I__289\ : InMux
    port map (
            O => \N__2385\,
            I => \N__2382\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2382\,
            I => \N__2379\
        );

    \I__287\ : Odrv4
    port map (
            O => \N__2379\,
            I => i2c_cmd_1_4
        );

    \I__286\ : InMux
    port map (
            O => \N__2376\,
            I => \N__2373\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2373\,
            I => \N__2370\
        );

    \I__284\ : Odrv4
    port map (
            O => \N__2370\,
            I => i2c_cmd_1_3
        );

    \I__283\ : InMux
    port map (
            O => \N__2367\,
            I => \bfn_1_4_0_\
        );

    \I__282\ : InMux
    port map (
            O => \N__2364\,
            I => \N__2360\
        );

    \I__281\ : InMux
    port map (
            O => \N__2363\,
            I => \N__2357\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2360\,
            I => \N__2352\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2357\,
            I => \N__2352\
        );

    \I__278\ : DummyBuf
    port map (
            O => \N__2352\,
            I => \hard0_SBDATo_0\
        );

    \I__277\ : InMux
    port map (
            O => \N__2349\,
            I => \N__2345\
        );

    \I__276\ : InMux
    port map (
            O => \N__2348\,
            I => \N__2342\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2345\,
            I => \N__2337\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2342\,
            I => \N__2337\
        );

    \I__273\ : DummyBuf
    port map (
            O => \N__2337\,
            I => \hard0_SBDATo_1\
        );

    \I__272\ : InMux
    port map (
            O => \N__2334\,
            I => \N__2330\
        );

    \I__271\ : InMux
    port map (
            O => \N__2333\,
            I => \N__2327\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2330\,
            I => \N__2322\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__2327\,
            I => \N__2322\
        );

    \I__268\ : DummyBuf
    port map (
            O => \N__2322\,
            I => \hard0_SBDATo_3\
        );

    \I__267\ : InMux
    port map (
            O => \N__2319\,
            I => \N__2315\
        );

    \I__266\ : InMux
    port map (
            O => \N__2318\,
            I => \N__2312\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2315\,
            I => \N__2307\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2312\,
            I => \N__2307\
        );

    \I__263\ : DummyBuf
    port map (
            O => \N__2307\,
            I => \hard0_SBDATo_4\
        );

    \I__262\ : InMux
    port map (
            O => \N__2304\,
            I => \N__2300\
        );

    \I__261\ : InMux
    port map (
            O => \N__2303\,
            I => \N__2297\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2300\,
            I => \N__2292\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__2297\,
            I => \N__2292\
        );

    \I__258\ : DummyBuf
    port map (
            O => \N__2292\,
            I => \hard0_SBDATo_5\
        );

    \I__257\ : InMux
    port map (
            O => \N__2289\,
            I => \N__2285\
        );

    \I__256\ : InMux
    port map (
            O => \N__2288\,
            I => \N__2282\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2285\,
            I => \N__2277\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2282\,
            I => \N__2277\
        );

    \I__253\ : DummyBuf
    port map (
            O => \N__2277\,
            I => \hard0_SBDATo_7\
        );

    \I__252\ : DummyBuf
    port map (
            O => \N__2274\,
            I => \N__2271\
        );

    \I__251\ : InMux
    port map (
            O => \N__2271\,
            I => \N__2268\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2268\,
            I => \N__2265\
        );

    \I__249\ : Odrv12
    port map (
            O => \N__2265\,
            I => \PWM_G\
        );

    \I__248\ : DummyBuf
    port map (
            O => \N__2262\,
            I => \N__2259\
        );

    \I__247\ : InMux
    port map (
            O => \N__2259\,
            I => \N__2256\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__2256\,
            I => \N__2253\
        );

    \I__245\ : Odrv12
    port map (
            O => \N__2253\,
            I => \PWM_R\
        );

    \I__244\ : CEMux
    port map (
            O => \N__2250\,
            I => \N__2247\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__2247\,
            I => \N__2243\
        );

    \I__242\ : CEMux
    port map (
            O => \N__2246\,
            I => \N__2240\
        );

    \I__241\ : Span4Mux_s1_h
    port map (
            O => \N__2243\,
            I => \N__2237\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__2240\,
            I => \N__2234\
        );

    \I__239\ : Span4Mux_h
    port map (
            O => \N__2237\,
            I => \N__2231\
        );

    \I__238\ : Odrv4
    port map (
            O => \N__2234\,
            I => n1815
        );

    \I__237\ : Odrv4
    port map (
            O => \N__2231\,
            I => n1815
        );

    \I__236\ : SRMux
    port map (
            O => \N__2226\,
            I => \N__2223\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__2223\,
            I => n1_adj_12
        );

    \I__234\ : DummyBuf
    port map (
            O => \N__2220\,
            I => \N__2217\
        );

    \I__233\ : InMux
    port map (
            O => \N__2217\,
            I => \N__2214\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__2214\,
            I => \N__2207\
        );

    \I__231\ : DummyBuf
    port map (
            O => \N__2213\,
            I => \N__2204\
        );

    \I__230\ : DummyBuf
    port map (
            O => \N__2212\,
            I => \N__2201\
        );

    \I__229\ : DummyBuf
    port map (
            O => \N__2211\,
            I => \N__2198\
        );

    \I__228\ : DummyBuf
    port map (
            O => \N__2210\,
            I => \N__2195\
        );

    \I__227\ : Span4Mux_s1_h
    port map (
            O => \N__2207\,
            I => \N__2192\
        );

    \I__226\ : InMux
    port map (
            O => \N__2204\,
            I => \N__2189\
        );

    \I__225\ : InMux
    port map (
            O => \N__2201\,
            I => \N__2186\
        );

    \I__224\ : InMux
    port map (
            O => \N__2198\,
            I => \N__2183\
        );

    \I__223\ : InMux
    port map (
            O => \N__2195\,
            I => \N__2180\
        );

    \I__222\ : Sp12to4
    port map (
            O => \N__2192\,
            I => \N__2177\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__2189\,
            I => \N__2168\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__2186\,
            I => \N__2168\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__2183\,
            I => \N__2168\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__2180\,
            I => \N__2168\
        );

    \I__217\ : Span12Mux_s8_v
    port map (
            O => \N__2177\,
            I => \N__2165\
        );

    \I__216\ : Sp12to4
    port map (
            O => \N__2168\,
            I => \N__2162\
        );

    \I__215\ : Span12Mux_h
    port map (
            O => \N__2165\,
            I => \N__2159\
        );

    \I__214\ : Odrv12
    port map (
            O => \N__2162\,
            I => \CONSTANT_ONE_NET\
        );

    \I__213\ : Odrv12
    port map (
            O => \N__2159\,
            I => \CONSTANT_ONE_NET\
        );

    \I__212\ : InMux
    port map (
            O => \N__2154\,
            I => \N__2151\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__2151\,
            I => n2967
        );

    \I__210\ : InMux
    port map (
            O => \N__2148\,
            I => \N__2145\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__2145\,
            I => n2966
        );

    \I__208\ : CascadeMux
    port map (
            O => \N__2142\,
            I => \n2811_cascade_\
        );

    \I__207\ : CascadeMux
    port map (
            O => \N__2139\,
            I => \n2821_cascade_\
        );

    \I__206\ : CascadeMux
    port map (
            O => \N__2136\,
            I => \n1_adj_12_cascade_\
        );

    \I__205\ : DummyBuf
    port map (
            O => \N__2133\,
            I => \N__2130\
        );

    \I__204\ : InMux
    port map (
            O => \N__2130\,
            I => \N__2127\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__2127\,
            I => \N__2124\
        );

    \I__202\ : Span12Mux_s3_v
    port map (
            O => \N__2124\,
            I => \N__2121\
        );

    \I__201\ : Odrv12
    port map (
            O => \N__2121\,
            I => \PWM_B\
        );

    \I__200\ : DummyBuf
    port map (
            O => \N__2118\,
            I => \N__2115\
        );

    \I__199\ : InMux
    port map (
            O => \N__2115\,
            I => \N__2112\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__2112\,
            I => \N__2109\
        );

    \I__197\ : Span12Mux_s10_h
    port map (
            O => \N__2109\,
            I => \N__2106\
        );

    \I__196\ : Span12Mux_v
    port map (
            O => \N__2106\,
            I => \N__2103\
        );

    \I__195\ : Odrv12
    port map (
            O => \N__2103\,
            I => sdain_i
        );

    \I__194\ : DummyBuf
    port map (
            O => \N__2100\,
            I => \N__2097\
        );

    \I__193\ : InMux
    port map (
            O => \N__2097\,
            I => \N__2094\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__2094\,
            I => \N__2091\
        );

    \I__191\ : Span4Mux_s2_v
    port map (
            O => \N__2091\,
            I => \N__2088\
        );

    \I__190\ : Sp12to4
    port map (
            O => \N__2088\,
            I => \N__2085\
        );

    \I__189\ : Span12Mux_s10_h
    port map (
            O => \N__2085\,
            I => \N__2082\
        );

    \I__188\ : Odrv12
    port map (
            O => \N__2082\,
            I => sclin_i
        );

    \I__187\ : CascadeMux
    port map (
            O => \N__2079\,
            I => \n2965_cascade_\
        );

    \I__186\ : CascadeMux
    port map (
            O => \N__2076\,
            I => \n2870_cascade_\
        );

    \I__185\ : CascadeMux
    port map (
            O => \N__2073\,
            I => \n6_adj_16_cascade_\
        );

    \I__184\ : IoInMux
    port map (
            O => \N__2070\,
            I => \N__2067\
        );

    \I__183\ : LocalMux
    port map (
            O => \N__2067\,
            I => \N__2064\
        );

    \I__182\ : IoSpan4Mux
    port map (
            O => \N__2064\,
            I => \N__2061\
        );

    \I__181\ : IoSpan4Mux
    port map (
            O => \N__2061\,
            I => \N__2058\
        );

    \I__180\ : Span4Mux_s3_v
    port map (
            O => \N__2058\,
            I => \N__2055\
        );

    \I__179\ : Sp12to4
    port map (
            O => \N__2055\,
            I => \N__2052\
        );

    \I__178\ : Odrv12
    port map (
            O => \N__2052\,
            I => \N__2049\
        );

    \I__177\ : DummyBuf
    port map (
            O => \N__2049\,
            I => sdaoe_i
        );

    \I__176\ : IoInMux
    port map (
            O => \N__2046\,
            I => \N__2043\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__2043\,
            I => \N__2040\
        );

    \I__174\ : IoSpan4Mux
    port map (
            O => \N__2040\,
            I => \N__2037\
        );

    \I__173\ : IoSpan4Mux
    port map (
            O => \N__2037\,
            I => \N__2034\
        );

    \I__172\ : Sp12to4
    port map (
            O => \N__2034\,
            I => \N__2031\
        );

    \I__171\ : Span12Mux_s5_v
    port map (
            O => \N__2031\,
            I => \N__2028\
        );

    \I__170\ : Odrv12
    port map (
            O => \N__2028\,
            I => \N__2025\
        );

    \I__169\ : DummyBuf
    port map (
            O => \N__2025\,
            I => sdaout_i
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2528,
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_4_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b00"
        )
    port map (
            CLKHFPU => \N__2212\,
            CLKHFEN => \N__2211\,
            CLKHF => n2981
        );

    \RGB_DRV\ : SB_RGBA_DRV
    generic map (
            RGB0_CURRENT => "0b000111",
            CURRENT_MODE => "0b0",
            RGB2_CURRENT => "0b000111",
            RGB1_CURRENT => "0b000111"
        )
    port map (
            RGBLEDEN => \N__2210\,
            RGB2PWM => \N__2133\,
            RGB1 => \LED_G_wire\,
            CURREN => \N__2220\,
            RGB2 => \LED_B_wire\,
            RGB1PWM => \N__2274\,
            RGB0PWM => \N__2262\,
            RGB0 => \LED_R_wire\
        );

    \I2C_1\ : SB_I2C_FIFO
    generic map (
            I2C_SLAVE_ADDR => "0b1000001"
        )
    port map (
            MRDCMPL => OPEN,
            DATO4 => \hard0_SBDATo_4\,
            WEI => \N__3564\,
            DATI3 => '0',
            TXFIFOAEMPTY => OPEN,
            DATO6 => \hard0_SBDATo_6\,
            DATO1 => \hard0_SBDATo_1\,
            DATI1 => '0',
            SDAOE => sdaoe_i,
            SDAI => \N__2118\,
            SCLOE => OPEN,
            DATO8 => OPEN,
            DATO0 => \hard0_SBDATo_0\,
            DATI8 => '0',
            DATI0 => '0',
            ADRI2 => \N__3522\,
            TXFIFOFULL => OPEN,
            TXFIFOEMPTY => OPEN,
            STBI => \N__3765\,
            RXFIFOFULL => OPEN,
            DATO3 => \hard0_SBDATo_3\,
            DATI7 => \N__3804\,
            ADRI1 => \N__3840\,
            ACKO => \hard0_SBACKo\,
            SDAO => sdaout_i,
            I2CWKUP => OPEN,
            I2CIRQ => OPEN,
            DATO2 => \hard0_SBDATo_2\,
            DATI6 => '0',
            CLKI => \N__3596\,
            ADRI0 => \N__3546\,
            RXFIFOAFULL => OPEN,
            FIFORST => '0',
            DATO5 => \hard0_SBDATo_5\,
            DATI5 => '0',
            SCLI => \N__2100\,
            DATI4 => \N__3687\,
            DATO7 => \hard0_SBDATo_7\,
            SCLO => OPEN,
            DATI2 => \N__3657\,
            SRWO => OPEN,
            RXFIFOEMPTY => OPEN,
            DATO9 => OPEN,
            DATI9 => '0',
            CSI => \N__2213\,
            ADRI3 => \N__3621\
        );

    \sysclk_GB\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3579\,
            GLOBALBUFFEROUTPUT => sysclk
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PWM_cnt_7__I_0_i9_2_lut_rep_47_LC_0_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2700\,
            in2 => \_gnd_net_\,
            in3 => \N__2719\,
            lcout => OPEN,
            ltout => \n2965_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1882_4_lut_LC_0_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001001"
        )
    port map (
            in0 => \N__2777\,
            in1 => \N__2421\,
            in2 => \N__2079\,
            in3 => \N__2154\,
            lcout => OPEN,
            ltout => \n2870_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1893_4_lut_LC_0_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2148\,
            in1 => \N__3015\,
            in2 => \N__2076\,
            in3 => \N__3384\,
            lcout => n2881,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_cnt_7__I_0_i6_3_lut_3_lut_LC_0_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__2735\,
            in1 => \_gnd_net_\,
            in2 => \N__2760\,
            in3 => \N__2420\,
            lcout => OPEN,
            ltout => \n6_adj_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_cnt_7__I_0_i8_3_lut_3_lut_LC_0_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2720\,
            in2 => \N__2073\,
            in3 => \N__2701\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_cnt_7__I_0_i4_4_lut_4_lut_LC_0_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001110"
        )
    port map (
            in0 => \N__2994\,
            in1 => \N__2940\,
            in2 => \N__2963\,
            in3 => \N__2981\,
            lcout => n4_adj_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_8_i7_2_lut_rep_49_LC_0_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2734\,
            in2 => \_gnd_net_\,
            in3 => \N__2754\,
            lcout => n2967,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_cnt_7__I_0_i11_2_lut_rep_48_LC_0_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3032\,
            in2 => \_gnd_net_\,
            in3 => \N__2876\,
            lcout => n2966,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \drv_cnt_i0_i1_LC_0_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001100110"
        )
    port map (
            in0 => \N__2580\,
            in1 => \N__2543\,
            in2 => \_gnd_net_\,
            in3 => \N__2514\,
            lcout => drv_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4256\,
            ce => \N__2598\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_11_LC_0_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3346\,
            in1 => \N__3145\,
            in2 => \_gnd_net_\,
            in3 => \N__3127\,
            lcout => OPEN,
            ltout => \n2811_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_6_LC_0_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__3364\,
            in1 => \N__3295\,
            in2 => \N__2142\,
            in3 => \N__3272\,
            lcout => OPEN,
            ltout => \n2821_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1846_4_lut_LC_0_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__3210\,
            in1 => \N__3313\,
            in2 => \N__2139\,
            in3 => \N__3184\,
            lcout => n105,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_0_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2672\,
            in2 => \_gnd_net_\,
            in3 => \N__2657\,
            lcout => n2819,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1926_2_lut_LC_0_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__3258\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3461\,
            lcout => n1_adj_12,
            ltout => \n1_adj_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_B_142_LC_0_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__2574\,
            in1 => \N__2551\,
            in2 => \N__2136\,
            in3 => \N__2515\,
            lcout => \PWM_B\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4258\,
            ce => \N__2250\,
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_8_LC_0_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__3460\,
            in1 => \N__3257\,
            in2 => \_gnd_net_\,
            in3 => \N__2615\,
            lcout => n1815,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_G_143_LC_0_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111001100"
        )
    port map (
            in0 => \N__2552\,
            in1 => \N__2584\,
            in2 => \_gnd_net_\,
            in3 => \N__2516\,
            lcout => \PWM_G\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4260\,
            ce => \N__2246\,
            sr => \N__2226\
        );

    \PWM_R_144_LC_0_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111110000"
        )
    port map (
            in0 => \N__2517\,
            in1 => \_gnd_net_\,
            in2 => \N__2589\,
            in3 => \N__2553\,
            lcout => \PWM_R\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4260\,
            ce => \N__2246\,
            sr => \N__2226\
        );

    \CONSTANT_ONE_LUT4_LC_0_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i10_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2348\,
            lcout => i2c_cmd_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4248\,
            ce => \N__4353\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i11_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4156\,
            lcout => i2c_cmd_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4248\,
            ce => \N__4353\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i12_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2333\,
            lcout => i2c_cmd_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4248\,
            ce => \N__4353\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i13_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2318\,
            lcout => i2c_cmd_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4248\,
            ce => \N__4353\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i14_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2303\,
            lcout => i2c_cmd_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4248\,
            ce => \N__4353\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i15_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4009\,
            lcout => i2c_cmd_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4248\,
            ce => \N__4353\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i16_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2288\,
            lcout => i2c_cmd_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4248\,
            ce => \N__4353\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i9_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2363\,
            lcout => i2c_cmd_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4248\,
            ce => \N__4353\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i1_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2364\,
            lcout => i2c_cmd_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4251\,
            ce => \N__3885\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i2_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2349\,
            lcout => i2c_cmd_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4251\,
            ce => \N__3885\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i4_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2334\,
            lcout => i2c_cmd_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4251\,
            ce => \N__3885\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i5_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2319\,
            lcout => i2c_cmd_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4251\,
            ce => \N__3885\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i6_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2304\,
            lcout => i2c_cmd_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4251\,
            ce => \N__3885\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i7_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4010\,
            lcout => i2c_cmd_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4251\,
            ce => \N__3885\,
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i8_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2289\,
            lcout => i2c_cmd_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4251\,
            ce => \N__3885\,
            sr => \_gnd_net_\
        );

    \PWM_duty_i0_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2448\,
            lcout => \PWM_duty_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4253\,
            ce => \N__3042\,
            sr => \_gnd_net_\
        );

    \PWM_duty_i1_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2439\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWM_duty_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4253\,
            ce => \N__3042\,
            sr => \_gnd_net_\
        );

    \PWM_duty_i2_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2430\,
            lcout => \PWM_duty_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4253\,
            ce => \N__3042\,
            sr => \_gnd_net_\
        );

    \PWM_duty_i5_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2412\,
            lcout => \PWM_duty_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4253\,
            ce => \N__3042\,
            sr => \_gnd_net_\
        );

    \PWM_duty_i6_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2403\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWM_duty_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4253\,
            ce => \N__3042\,
            sr => \_gnd_net_\
        );

    \PWM_duty_i7_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2394\,
            lcout => \PWM_duty_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4253\,
            ce => \N__3042\,
            sr => \_gnd_net_\
        );

    \PWM_duty_i4_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2385\,
            lcout => \PWM_duty_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4253\,
            ce => \N__3042\,
            sr => \_gnd_net_\
        );

    \PWM_duty_i3_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2376\,
            lcout => \PWM_duty_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4253\,
            ce => \N__3042\,
            sr => \_gnd_net_\
        );

    \PWM_cnt__i0_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2962\,
            in2 => \_gnd_net_\,
            in3 => \N__2367\,
            lcout => \PWM_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_1_4_0_\,
            carryout => n2514,
            clk => \N__4254\,
            ce => \N__2457\,
            sr => \N__3435\
        );

    \PWM_cnt__i1_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2982\,
            in2 => \_gnd_net_\,
            in3 => \N__2478\,
            lcout => \PWM_cnt_1\,
            ltout => OPEN,
            carryin => n2514,
            carryout => n2515,
            clk => \N__4254\,
            ce => \N__2457\,
            sr => \N__3435\
        );

    \PWM_cnt__i2_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2778\,
            in2 => \_gnd_net_\,
            in3 => \N__2475\,
            lcout => \PWM_cnt_2\,
            ltout => OPEN,
            carryin => n2515,
            carryout => n2516,
            clk => \N__4254\,
            ce => \N__2457\,
            sr => \N__3435\
        );

    \PWM_cnt__i3_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2759\,
            in2 => \_gnd_net_\,
            in3 => \N__2472\,
            lcout => \PWM_cnt_3\,
            ltout => OPEN,
            carryin => n2516,
            carryout => n2517,
            clk => \N__4254\,
            ce => \N__2457\,
            sr => \N__3435\
        );

    \PWM_cnt__i4_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2703\,
            in2 => \_gnd_net_\,
            in3 => \N__2469\,
            lcout => \PWM_cnt_4\,
            ltout => OPEN,
            carryin => n2517,
            carryout => n2518,
            clk => \N__4254\,
            ce => \N__2457\,
            sr => \N__3435\
        );

    \PWM_cnt__i5_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2877\,
            in2 => \_gnd_net_\,
            in3 => \N__2466\,
            lcout => \PWM_cnt_5\,
            ltout => OPEN,
            carryin => n2518,
            carryout => n2519,
            clk => \N__4254\,
            ce => \N__2457\,
            sr => \N__3435\
        );

    \PWM_cnt__i6_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2901\,
            in2 => \_gnd_net_\,
            in3 => \N__2463\,
            lcout => \PWM_cnt_6\,
            ltout => OPEN,
            carryin => n2519,
            carryout => n2520,
            clk => \N__4254\,
            ce => \N__2457\,
            sr => \N__3435\
        );

    \PWM_cnt__i7_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3408\,
            in2 => \_gnd_net_\,
            in3 => \N__2460\,
            lcout => \PWM_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4254\,
            ce => \N__2457\,
            sr => \N__3435\
        );

    \i1921_2_lut_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__3463\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3260\,
            lcout => n1831,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \drv_cnt_i0_i0_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001101100"
        )
    port map (
            in0 => \N__3261\,
            in1 => \N__2545\,
            in2 => \N__2616\,
            in3 => \N__3464\,
            lcout => drv_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4255\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_cnt_7__I_0_i12_3_lut_3_lut_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3407\,
            in2 => \N__2793\,
            in3 => \N__3426\,
            lcout => OPEN,
            ltout => \n12_adj_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_cnt_7__I_0_i14_3_lut_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3003\,
            in2 => \N__2634\,
            in3 => \N__2631\,
            lcout => OPEN,
            ltout => \n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1049_3_lut_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2625\,
            in2 => \N__2619\,
            in3 => \N__3488\,
            lcout => n2012,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_8_i13_2_lut_rep_50_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2922\,
            in2 => \_gnd_net_\,
            in3 => \N__2898\,
            lcout => n2968,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_rep_37_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__3462\,
            in1 => \N__3259\,
            in2 => \_gnd_net_\,
            in3 => \N__2611\,
            lcout => n2955,
            ltout => \n2955_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \drv_cnt_i0_i2_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110000000"
        )
    port map (
            in0 => \N__2588\,
            in1 => \N__2544\,
            in2 => \N__2520\,
            in3 => \N__2508\,
            lcout => drv_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4255\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \drv_clk_counter_526__i0_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3329\,
            in2 => \_gnd_net_\,
            in3 => \N__2487\,
            lcout => drv_clk_counter_0,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => n2521,
            clk => \N__4257\,
            ce => 'H',
            sr => \N__3164\
        );

    \drv_clk_counter_526__i1_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3348\,
            in2 => \_gnd_net_\,
            in3 => \N__2484\,
            lcout => drv_clk_counter_1,
            ltout => OPEN,
            carryin => n2521,
            carryout => n2522,
            clk => \N__4257\,
            ce => 'H',
            sr => \N__3164\
        );

    \drv_clk_counter_526__i2_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3147\,
            in2 => \_gnd_net_\,
            in3 => \N__2481\,
            lcout => drv_clk_counter_2,
            ltout => OPEN,
            carryin => n2522,
            carryout => n2523,
            clk => \N__4257\,
            ce => 'H',
            sr => \N__3164\
        );

    \drv_clk_counter_526__i3_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3129\,
            in2 => \_gnd_net_\,
            in3 => \N__2682\,
            lcout => drv_clk_counter_3,
            ltout => OPEN,
            carryin => n2523,
            carryout => n2524,
            clk => \N__4257\,
            ce => 'H',
            sr => \N__3164\
        );

    \drv_clk_counter_526__i4_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3366\,
            in2 => \_gnd_net_\,
            in3 => \N__2679\,
            lcout => drv_clk_counter_4,
            ltout => OPEN,
            carryin => n2524,
            carryout => n2525,
            clk => \N__4257\,
            ce => 'H',
            sr => \N__3164\
        );

    \drv_clk_counter_526__i5_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3297\,
            in2 => \_gnd_net_\,
            in3 => \N__2676\,
            lcout => drv_clk_counter_5,
            ltout => OPEN,
            carryin => n2525,
            carryout => n2526,
            clk => \N__4257\,
            ce => 'H',
            sr => \N__3164\
        );

    \drv_clk_counter_526__i6_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2673\,
            in2 => \_gnd_net_\,
            in3 => \N__2661\,
            lcout => drv_clk_counter_6,
            ltout => OPEN,
            carryin => n2526,
            carryout => n2527,
            clk => \N__4257\,
            ce => 'H',
            sr => \N__3164\
        );

    \drv_clk_counter_526__i7_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2658\,
            in2 => \_gnd_net_\,
            in3 => \N__2646\,
            lcout => drv_clk_counter_7,
            ltout => OPEN,
            carryin => n2527,
            carryout => n2528,
            clk => \N__4257\,
            ce => 'H',
            sr => \N__3164\
        );

    \drv_clk_counter_526__i8_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3315\,
            in2 => \_gnd_net_\,
            in3 => \N__2643\,
            lcout => drv_clk_counter_8,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => n2529,
            clk => \N__4259\,
            ce => 'H',
            sr => \N__3168\
        );

    \drv_clk_counter_526__i9_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3186\,
            in2 => \_gnd_net_\,
            in3 => \N__2640\,
            lcout => drv_clk_counter_9,
            ltout => OPEN,
            carryin => n2529,
            carryout => n2530,
            clk => \N__4259\,
            ce => 'H',
            sr => \N__3168\
        );

    \drv_clk_counter_526__i10_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3209\,
            in2 => \_gnd_net_\,
            in3 => \N__2637\,
            lcout => drv_clk_counter_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4259\,
            ce => 'H',
            sr => \N__3168\
        );

    \i1852_2_lut_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2822\,
            in2 => \_gnd_net_\,
            in3 => \N__2810\,
            lcout => OPEN,
            ltout => \n2838_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1871_4_lut_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2835\,
            in1 => \N__2844\,
            in2 => \N__2847\,
            in3 => \N__2802\,
            lcout => n2858,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_21_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2843\,
            in2 => \_gnd_net_\,
            in3 => \N__2801\,
            lcout => OPEN,
            ltout => \n6_adj_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2834\,
            in1 => \N__2823\,
            in2 => \N__2814\,
            in3 => \N__2811\,
            lcout => n2247,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2c_cmd_0___i3_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4160\,
            lcout => i2c_cmd_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4249\,
            ce => \N__3881\,
            sr => \_gnd_net_\
        );

    \PWM_cnt_7__I_0_i10_3_lut_3_lut_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__2899\,
            in1 => \N__2920\,
            in2 => \_gnd_net_\,
            in3 => \N__3031\,
            lcout => n10_adj_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i30_4_lut_3_lut_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101100110"
        )
    port map (
            in0 => \N__3058\,
            in1 => \N__3091\,
            in2 => \_gnd_net_\,
            in3 => \N__3077\,
            lcout => OPEN,
            ltout => \n17_adj_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cmd_decoded_156_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__3105\,
            in1 => \N__4073\,
            in2 => \N__2781\,
            in3 => \N__4338\,
            lcout => cmd_decoded,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4252\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_8_i6_3_lut_3_lut_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__2776\,
            in1 => \N__2758\,
            in2 => \_gnd_net_\,
            in3 => \N__2736\,
            lcout => OPEN,
            ltout => \n6_adj_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_8_i8_3_lut_3_lut_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2721\,
            in2 => \N__2706\,
            in3 => \N__2702\,
            lcout => n8_adj_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1286_2_lut_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3076\,
            in2 => \_gnd_net_\,
            in3 => \N__3104\,
            lcout => OPEN,
            ltout => \n2250_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \motor_on_158_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110100010"
        )
    port map (
            in0 => \N__3243\,
            in1 => \N__3062\,
            in2 => \N__3096\,
            in3 => \N__3093\,
            lcout => motor_on,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4252\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__3092\,
            in1 => \N__3078\,
            in2 => \N__3063\,
            in3 => \N__3048\,
            lcout => n1778,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1895_3_lut_3_lut_4_lut_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001001"
        )
    port map (
            in0 => \N__2875\,
            in1 => \N__3033\,
            in2 => \N__3383\,
            in3 => \N__3014\,
            lcout => n2883,
            ltout => \n2883_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_8_i14_3_lut_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2928\,
            in2 => \N__2997\,
            in3 => \N__2853\,
            lcout => n14_adj_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_8_i4_4_lut_4_lut_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011011100"
        )
    port map (
            in0 => \N__2993\,
            in1 => \N__2980\,
            in2 => \N__2964\,
            in3 => \N__2939\,
            lcout => n4_adj_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_8_i10_3_lut_3_lut_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__2921\,
            in1 => \N__2900\,
            in2 => \_gnd_net_\,
            in3 => \N__2874\,
            lcout => OPEN,
            ltout => \n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_8_i12_3_lut_3_lut_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101010000"
        )
    port map (
            in0 => \N__3422\,
            in1 => \_gnd_net_\,
            in2 => \N__2856\,
            in3 => \N__3406\,
            lcout => n12_adj_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_8_i16_3_lut_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3498\,
            in1 => \N__3492\,
            in2 => \_gnd_net_\,
            in3 => \N__3477\,
            lcout => OPEN,
            ltout => \n104_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_20_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3242\,
            in2 => \N__3471\,
            in3 => \N__3468\,
            lcout => n1921,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_8_i15_2_lut_rep_51_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3421\,
            in2 => \_gnd_net_\,
            in3 => \N__3405\,
            lcout => n2969,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_9_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__3365\,
            in1 => \N__3347\,
            in2 => \N__3330\,
            in3 => \N__3111\,
            lcout => OPEN,
            ltout => \n2810_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_10_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__3314\,
            in1 => \N__3296\,
            in2 => \N__3279\,
            in3 => \N__3276\,
            lcout => OPEN,
            ltout => \n2820_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i248_4_lut_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111010101"
        )
    port map (
            in0 => \N__3249\,
            in1 => \N__3208\,
            in2 => \N__3189\,
            in3 => \N__3185\,
            lcout => n953,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_rep_45_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3146\,
            in2 => \_gnd_net_\,
            in3 => \N__3128\,
            lcout => n2963,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_12_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__4703\,
            in1 => \N__4932\,
            in2 => \_gnd_net_\,
            in3 => \N__4482\,
            lcout => OPEN,
            ltout => \n2824_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \soft_SBADRi_i3_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111100101111"
        )
    port map (
            in0 => \N__3614\,
            in1 => \N__3734\,
            in2 => \N__3624\,
            in3 => \N__4484\,
            lcout => \hard_SBADRi_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_n2981_THRU_LUT4_0_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3600\,
            lcout => \GB_BUFFER_n2981_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i745_2_lut_rep_42_4_lut_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__4483\,
            in1 => \N__4830\,
            in2 => \N__4719\,
            in3 => \N__4596\,
            lcout => OPEN,
            ltout => \n2960_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \hard_SBWRi_147_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__4933\,
            in1 => \N__3560\,
            in2 => \N__3567\,
            in3 => \N__4707\,
            lcout => \hard_SBWRi\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \soft_SBADRi_i0_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__3630\,
            in1 => \N__3701\,
            in2 => \N__3545\,
            in3 => \N__3866\,
            lcout => \hard_SBADRi_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1256_2_lut_rep_53_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4700\,
            in2 => \_gnd_net_\,
            in3 => \N__4583\,
            lcout => n2971,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i28_4_lut_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010000"
        )
    port map (
            in0 => \N__4585\,
            in1 => \N__3865\,
            in2 => \N__3518\,
            in3 => \N__4832\,
            lcout => OPEN,
            ltout => \n12_adj_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \soft_SBADRi_i2_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__4481\,
            in1 => \N__3514\,
            in2 => \N__3525\,
            in3 => \N__4702\,
            lcout => \hard_SBADRi_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i29_3_lut_4_lut_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__4931\,
            in1 => \N__4478\,
            in2 => \N__3680\,
            in3 => \N__4831\,
            lcout => OPEN,
            ltout => \n13_adj_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \hard_SBDATi_i4_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__4480\,
            in1 => \N__3702\,
            in2 => \N__3690\,
            in3 => \N__3676\,
            lcout => \hard_SBDATi_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i28_4_lut_4_lut_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001010000"
        )
    port map (
            in0 => \N__4584\,
            in1 => \N__3864\,
            in2 => \N__3650\,
            in3 => \N__4833\,
            lcout => OPEN,
            ltout => \n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \hard_SBDATi_i2_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__4479\,
            in1 => \N__3646\,
            in2 => \N__3660\,
            in3 => \N__4701\,
            lcout => \hard_SBDATi_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1923_2_lut_rep_41_4_lut_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4426\,
            in1 => \N__4815\,
            in2 => \N__4716\,
            in3 => \N__4594\,
            lcout => n2959,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__4425\,
            in1 => \N__4816\,
            in2 => \N__4717\,
            in3 => \N__4595\,
            lcout => n15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1241_2_lut_rep_54_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4405\,
            in2 => \_gnd_net_\,
            in3 => \N__4879\,
            lcout => n2972,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2c_steps_i3_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__4051\,
            in1 => \N__4470\,
            in2 => \_gnd_net_\,
            in3 => \N__4841\,
            lcout => i2c_steps_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4250\,
            ce => 'H',
            sr => \N__3924\
        );

    \i2c_cnt_523_524__i2_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011110000"
        )
    port map (
            in0 => \N__3944\,
            in1 => \_gnd_net_\,
            in2 => \N__3966\,
            in3 => \N__3894\,
            lcout => i2c_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_587_i3_2_lut_rep_56_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3960\,
            in2 => \_gnd_net_\,
            in3 => \N__3942\,
            lcout => OPEN,
            ltout => \n2974_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i36_4_lut_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100001100"
        )
    port map (
            in0 => \N__4808\,
            in1 => \N__4550\,
            in2 => \N__3771\,
            in3 => \N__3981\,
            lcout => n31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2c_cnt_523_524__i1_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100100010"
        )
    port map (
            in0 => \N__3893\,
            in1 => \N__3961\,
            in2 => \_gnd_net_\,
            in3 => \N__3943\,
            lcout => i2c_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1279_2_lut_3_lut_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4809\,
            in1 => \N__4671\,
            in2 => \_gnd_net_\,
            in3 => \N__4552\,
            lcout => n2243,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_rep_52_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4810\,
            in1 => \N__4672\,
            in2 => \_gnd_net_\,
            in3 => \N__4551\,
            lcout => n2970,
            ltout => \n2970_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \hard_SBSTBi_148_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111010"
        )
    port map (
            in0 => \N__3761\,
            in1 => \N__4934\,
            in2 => \N__3768\,
            in3 => \N__4471\,
            lcout => \hard_SBSTBi\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_13_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__4930\,
            in1 => \N__3708\,
            in2 => \N__4718\,
            in3 => \N__3747\,
            lcout => OPEN,
            ltout => \n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110011"
        )
    port map (
            in0 => \N__3741\,
            in1 => \N__3735\,
            in2 => \N__3720\,
            in3 => \N__4475\,
            lcout => n1887,
            ltout => \n1887_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2c_steps_i2_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011110011101100"
        )
    port map (
            in0 => \N__3920\,
            in1 => \N__4708\,
            in2 => \N__3717\,
            in3 => \N__3714\,
            lcout => i2c_steps_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1240_2_lut_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4554\,
            in1 => \_gnd_net_\,
            in2 => \N__4834\,
            in3 => \_gnd_net_\,
            lcout => n1852,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__4959\,
            in1 => \N__4799\,
            in2 => \_gnd_net_\,
            in3 => \N__4553\,
            lcout => n22_adj_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2c_steps_i1_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111011110000"
        )
    port map (
            in0 => \N__4555\,
            in1 => \N__3919\,
            in2 => \N__4835\,
            in3 => \N__3900\,
            lcout => i2c_steps_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_17_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__4476\,
            in1 => \N__4052\,
            in2 => \_gnd_net_\,
            in3 => \N__4800\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4801\,
            in1 => \N__4941\,
            in2 => \N__4056\,
            in3 => \N__4477\,
            lcout => n1779,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i29_4_lut_4_lut_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001010000"
        )
    port map (
            in0 => \N__4827\,
            in1 => \N__3867\,
            in2 => \N__3830\,
            in3 => \N__4561\,
            lcout => OPEN,
            ltout => \n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_14_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__3826\,
            in1 => \N__4670\,
            in2 => \N__3846\,
            in3 => \N__4409\,
            lcout => OPEN,
            ltout => \n4_adj_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \soft_SBADRi_i1_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__4023\,
            in1 => \N__4883\,
            in2 => \N__3843\,
            in3 => \N__4563\,
            lcout => \hard_SBADRi_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111011100"
        )
    port map (
            in0 => \N__4881\,
            in1 => \N__4406\,
            in2 => \N__4842\,
            in3 => \N__4669\,
            lcout => n4_adj_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i29_3_lut_4_lut_adj_1_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__4407\,
            in1 => \N__4882\,
            in2 => \N__3794\,
            in3 => \N__4562\,
            lcout => OPEN,
            ltout => \n13_adj_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \hard_SBDATi_i7_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__3790\,
            in1 => \N__4029\,
            in2 => \N__3807\,
            in3 => \N__4410\,
            lcout => \hard_SBDATi_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_rep_43_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4668\,
            in1 => \N__4880\,
            in2 => \_gnd_net_\,
            in3 => \N__4560\,
            lcout => n2961,
            ltout => \n2961_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_4_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4074\,
            in1 => \N__4408\,
            in2 => \N__4059\,
            in3 => \N__4826\,
            lcout => n2016,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_rep_38_3_lut_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__4424\,
            in1 => \N__4050\,
            in2 => \_gnd_net_\,
            in3 => \N__4839\,
            lcout => n2956,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1844_2_lut_rep_55_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4715\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4840\,
            lcout => n2973,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_rep_44_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4423\,
            in2 => \_gnd_net_\,
            in3 => \N__4714\,
            lcout => n2962,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_55_i7_3_lut_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3983\,
            in1 => \N__4017\,
            in2 => \_gnd_net_\,
            in3 => \N__4929\,
            lcout => OPEN,
            ltout => \i2c_stat_7_N_205_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2c_stat_i6_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__4086\,
            in1 => \N__4101\,
            in2 => \N__3987\,
            in3 => \N__3984\,
            lcout => i2c_stat_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4240\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1293_3_lut_4_lut_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__3982\,
            in1 => \N__3965\,
            in2 => \N__4582\,
            in3 => \N__3945\,
            lcout => n2534,
            ltout => \n2534_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i58_4_lut_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__4696\,
            in1 => \N__4960\,
            in2 => \N__3927\,
            in3 => \N__4825\,
            lcout => OPEN,
            ltout => \n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__4559\,
            in1 => \_gnd_net_\,
            in2 => \N__4164\,
            in3 => \N__4928\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_55_i3_3_lut_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4161\,
            in1 => \N__4926\,
            in2 => \_gnd_net_\,
            in3 => \N__4961\,
            lcout => \i2c_stat_7_N_205_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1863_4_lut_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__4580\,
            in1 => \N__4712\,
            in2 => \N__4935\,
            in3 => \N__4828\,
            lcout => n2850,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_7_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4710\,
            in1 => \N__4473\,
            in2 => \_gnd_net_\,
            in3 => \N__4579\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i60_3_lut_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4922\,
            in1 => \N__4134\,
            in2 => \_gnd_net_\,
            in3 => \N__4829\,
            lcout => OPEN,
            ltout => \n2840_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_2_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000000000"
        )
    port map (
            in0 => \N__4713\,
            in1 => \N__4128\,
            in2 => \N__4119\,
            in3 => \N__4581\,
            lcout => OPEN,
            ltout => \n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2c_steps_i0_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110001"
        )
    port map (
            in0 => \N__4474\,
            in1 => \N__4116\,
            in2 => \N__4110\,
            in3 => \N__4107\,
            lcout => i2c_steps_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4241\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_rep_40_3_lut_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__4711\,
            in1 => \N__4472\,
            in2 => \_gnd_net_\,
            in3 => \N__4578\,
            lcout => n2958,
            ltout => \n2958_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2c_stat_i2_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__4962\,
            in1 => \N__4095\,
            in2 => \N__4089\,
            in3 => \N__4085\,
            lcout => i2c_stat_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4241\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_rep_46_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4319\,
            in2 => \_gnd_net_\,
            in3 => \N__4294\,
            lcout => n2964,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_rep_39_4_lut_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4927\,
            in1 => \N__4811\,
            in2 => \N__4709\,
            in3 => \N__4564\,
            lcout => OPEN,
            ltout => \n2957_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_5_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4323\,
            in1 => \N__4296\,
            in2 => \N__4488\,
            in3 => \N__4485\,
            lcout => n1780,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__4295\,
            in1 => \_gnd_net_\,
            in2 => \N__4326\,
            in3 => \N__4275\,
            lcout => n1730,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2c_cmd_cnt_525__i1_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__4298\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4324\,
            lcout => i2c_cmd_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4245\,
            ce => \N__4191\,
            sr => \N__4176\
        );

    \i2c_cmd_cnt_525__i0_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4297\,
            lcout => i2c_cmd_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4245\,
            ce => \N__4191\,
            sr => \N__4176\
        );

    \i2c_cmd_cnt_525__i2_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__4325\,
            in1 => \N__4274\,
            in2 => \_gnd_net_\,
            in3 => \N__4299\,
            lcout => i2c_cmd_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4245\,
            ce => \N__4191\,
            sr => \N__4176\
        );
end \INTERFACE\;
